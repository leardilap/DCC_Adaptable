-- de2i_150_qsys.vhd

-- Generated using ACDS version 14.0 200 at 2015.10.12.22:26:00

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity de2i_150_qsys is
	port (
		clk_clk                                    : in  std_logic                     := '0';             --                        clk.clk
		reset_reset_n                              : in  std_logic                     := '0';             --                      reset.reset_n
		pcie_ip_reconfig_togxb_data                : in  std_logic_vector(3 downto 0)  := (others => '0'); --     pcie_ip_reconfig_togxb.data
		pcie_ip_refclk_export                      : in  std_logic                     := '0';             --             pcie_ip_refclk.export
		pcie_ip_test_in_test_in                    : in  std_logic_vector(39 downto 0) := (others => '0'); --            pcie_ip_test_in.test_in
		pcie_ip_pcie_rstn_export                   : in  std_logic                     := '0';             --          pcie_ip_pcie_rstn.export
		pcie_ip_clocks_sim_clk250_export           : out std_logic;                                        --         pcie_ip_clocks_sim.clk250_export
		pcie_ip_clocks_sim_clk500_export           : out std_logic;                                        --                           .clk500_export
		pcie_ip_clocks_sim_clk125_export           : out std_logic;                                        --                           .clk125_export
		pcie_ip_reconfig_busy_busy_altgxb_reconfig : in  std_logic                     := '0';             --      pcie_ip_reconfig_busy.busy_altgxb_reconfig
		pcie_ip_pipe_ext_pipe_mode                 : in  std_logic                     := '0';             --           pcie_ip_pipe_ext.pipe_mode
		pcie_ip_pipe_ext_phystatus_ext             : in  std_logic                     := '0';             --                           .phystatus_ext
		pcie_ip_pipe_ext_rate_ext                  : out std_logic;                                        --                           .rate_ext
		pcie_ip_pipe_ext_powerdown_ext             : out std_logic_vector(1 downto 0);                     --                           .powerdown_ext
		pcie_ip_pipe_ext_txdetectrx_ext            : out std_logic;                                        --                           .txdetectrx_ext
		pcie_ip_pipe_ext_rxelecidle0_ext           : in  std_logic                     := '0';             --                           .rxelecidle0_ext
		pcie_ip_pipe_ext_rxdata0_ext               : in  std_logic_vector(7 downto 0)  := (others => '0'); --                           .rxdata0_ext
		pcie_ip_pipe_ext_rxstatus0_ext             : in  std_logic_vector(2 downto 0)  := (others => '0'); --                           .rxstatus0_ext
		pcie_ip_pipe_ext_rxvalid0_ext              : in  std_logic                     := '0';             --                           .rxvalid0_ext
		pcie_ip_pipe_ext_rxdatak0_ext              : in  std_logic                     := '0';             --                           .rxdatak0_ext
		pcie_ip_pipe_ext_txdata0_ext               : out std_logic_vector(7 downto 0);                     --                           .txdata0_ext
		pcie_ip_pipe_ext_txdatak0_ext              : out std_logic;                                        --                           .txdatak0_ext
		pcie_ip_pipe_ext_rxpolarity0_ext           : out std_logic;                                        --                           .rxpolarity0_ext
		pcie_ip_pipe_ext_txcompl0_ext              : out std_logic;                                        --                           .txcompl0_ext
		pcie_ip_pipe_ext_txelecidle0_ext           : out std_logic;                                        --                           .txelecidle0_ext
		pcie_ip_rx_in_rx_datain_0                  : in  std_logic                     := '0';             --              pcie_ip_rx_in.rx_datain_0
		pcie_ip_tx_out_tx_dataout_0                : out std_logic;                                        --             pcie_ip_tx_out.tx_dataout_0
		pcie_ip_reconfig_fromgxb_0_data            : out std_logic_vector(4 downto 0);                     -- pcie_ip_reconfig_fromgxb_0.data
		led_external_connection_export             : out std_logic_vector(3 downto 0);                     --    led_external_connection.export
		button_external_connection_export          : in  std_logic_vector(3 downto 0)  := (others => '0'); -- button_external_connection.export
		fir_memory_s2_address                      : in  std_logic_vector(9 downto 0)  := (others => '0'); --              fir_memory_s2.address
		fir_memory_s2_chipselect                   : in  std_logic                     := '0';             --                           .chipselect
		fir_memory_s2_clken                        : in  std_logic                     := '0';             --                           .clken
		fir_memory_s2_write                        : in  std_logic                     := '0';             --                           .write
		fir_memory_s2_readdata                     : out std_logic_vector(31 downto 0);                    --                           .readdata
		fir_memory_s2_writedata                    : in  std_logic_vector(31 downto 0) := (others => '0'); --                           .writedata
		fir_memory_s2_byteenable                   : in  std_logic_vector(3 downto 0)  := (others => '0'); --                           .byteenable
		fir_memory_clk2_clk                        : in  std_logic                     := '0';             --            fir_memory_clk2.clk
		fir_memory_reset2_reset                    : in  std_logic                     := '0';             --          fir_memory_reset2.reset
		fir_memory_reset2_reset_req                : in  std_logic                     := '0';             --                           .reset_req
		interpo_4_0_s2_address                     : in  std_logic_vector(4 downto 0)  := (others => '0'); --             interpo_4_0_s2.address
		interpo_4_0_s2_chipselect                  : in  std_logic                     := '0';             --                           .chipselect
		interpo_4_0_s2_clken                       : in  std_logic                     := '0';             --                           .clken
		interpo_4_0_s2_write                       : in  std_logic                     := '0';             --                           .write
		interpo_4_0_s2_readdata                    : out std_logic_vector(31 downto 0);                    --                           .readdata
		interpo_4_0_s2_writedata                   : in  std_logic_vector(31 downto 0) := (others => '0'); --                           .writedata
		interpo_4_0_s2_byteenable                  : in  std_logic_vector(3 downto 0)  := (others => '0'); --                           .byteenable
		interpo_4_0_clk2_clk                       : in  std_logic                     := '0';             --           interpo_4_0_clk2.clk
		interpo_4_0_reset2_reset                   : in  std_logic                     := '0';             --         interpo_4_0_reset2.reset
		interpo_4_0_reset2_reset_req               : in  std_logic                     := '0';             --                           .reset_req
		interpo_5_0_s2_address                     : in  std_logic_vector(5 downto 0)  := (others => '0'); --             interpo_5_0_s2.address
		interpo_5_0_s2_chipselect                  : in  std_logic                     := '0';             --                           .chipselect
		interpo_5_0_s2_clken                       : in  std_logic                     := '0';             --                           .clken
		interpo_5_0_s2_write                       : in  std_logic                     := '0';             --                           .write
		interpo_5_0_s2_readdata                    : out std_logic_vector(31 downto 0);                    --                           .readdata
		interpo_5_0_s2_writedata                   : in  std_logic_vector(31 downto 0) := (others => '0'); --                           .writedata
		interpo_5_0_s2_byteenable                  : in  std_logic_vector(3 downto 0)  := (others => '0'); --                           .byteenable
		interpo_5_0_clk2_clk                       : in  std_logic                     := '0';             --           interpo_5_0_clk2.clk
		interpo_5_0_reset2_reset                   : in  std_logic                     := '0';             --         interpo_5_0_reset2.reset
		interpo_5_0_reset2_reset_req               : in  std_logic                     := '0';             --                           .reset_req
		interpo_5_1_clk2_clk                       : in  std_logic                     := '0';             --           interpo_5_1_clk2.clk
		interpo_5_1_s2_address                     : in  std_logic_vector(5 downto 0)  := (others => '0'); --             interpo_5_1_s2.address
		interpo_5_1_s2_chipselect                  : in  std_logic                     := '0';             --                           .chipselect
		interpo_5_1_s2_clken                       : in  std_logic                     := '0';             --                           .clken
		interpo_5_1_s2_write                       : in  std_logic                     := '0';             --                           .write
		interpo_5_1_s2_readdata                    : out std_logic_vector(31 downto 0);                    --                           .readdata
		interpo_5_1_s2_writedata                   : in  std_logic_vector(31 downto 0) := (others => '0'); --                           .writedata
		interpo_5_1_s2_byteenable                  : in  std_logic_vector(3 downto 0)  := (others => '0'); --                           .byteenable
		interpo_5_1_reset2_reset                   : in  std_logic                     := '0';             --         interpo_5_1_reset2.reset
		interpo_5_1_reset2_reset_req               : in  std_logic                     := '0';             --                           .reset_req
		interpo_5_2_s2_address                     : in  std_logic_vector(5 downto 0)  := (others => '0'); --             interpo_5_2_s2.address
		interpo_5_2_s2_chipselect                  : in  std_logic                     := '0';             --                           .chipselect
		interpo_5_2_s2_clken                       : in  std_logic                     := '0';             --                           .clken
		interpo_5_2_s2_write                       : in  std_logic                     := '0';             --                           .write
		interpo_5_2_s2_readdata                    : out std_logic_vector(31 downto 0);                    --                           .readdata
		interpo_5_2_s2_writedata                   : in  std_logic_vector(31 downto 0) := (others => '0'); --                           .writedata
		interpo_5_2_s2_byteenable                  : in  std_logic_vector(3 downto 0)  := (others => '0'); --                           .byteenable
		interpo_5_2_clk2_clk                       : in  std_logic                     := '0';             --           interpo_5_2_clk2.clk
		interpo_5_2_reset2_reset                   : in  std_logic                     := '0';             --         interpo_5_2_reset2.reset
		interpo_5_2_reset2_reset_req               : in  std_logic                     := '0';             --                           .reset_req
		interpo_5_3_s2_address                     : in  std_logic_vector(5 downto 0)  := (others => '0'); --             interpo_5_3_s2.address
		interpo_5_3_s2_chipselect                  : in  std_logic                     := '0';             --                           .chipselect
		interpo_5_3_s2_clken                       : in  std_logic                     := '0';             --                           .clken
		interpo_5_3_s2_write                       : in  std_logic                     := '0';             --                           .write
		interpo_5_3_s2_readdata                    : out std_logic_vector(31 downto 0);                    --                           .readdata
		interpo_5_3_s2_writedata                   : in  std_logic_vector(31 downto 0) := (others => '0'); --                           .writedata
		interpo_5_3_s2_byteenable                  : in  std_logic_vector(3 downto 0)  := (others => '0'); --                           .byteenable
		interpo_5_3_clk2_clk                       : in  std_logic                     := '0';             --           interpo_5_3_clk2.clk
		interpo_5_3_reset2_reset                   : in  std_logic                     := '0';             --         interpo_5_3_reset2.reset
		interpo_5_3_reset2_reset_req               : in  std_logic                     := '0';             --                           .reset_req
		adapt_fir_mem_s2_address                   : in  std_logic_vector(8 downto 0)  := (others => '0'); --           adapt_fir_mem_s2.address
		adapt_fir_mem_s2_chipselect                : in  std_logic                     := '0';             --                           .chipselect
		adapt_fir_mem_s2_clken                     : in  std_logic                     := '0';             --                           .clken
		adapt_fir_mem_s2_write                     : in  std_logic                     := '0';             --                           .write
		adapt_fir_mem_s2_readdata                  : out std_logic_vector(31 downto 0);                    --                           .readdata
		adapt_fir_mem_s2_writedata                 : in  std_logic_vector(31 downto 0) := (others => '0'); --                           .writedata
		adapt_fir_mem_s2_byteenable                : in  std_logic_vector(3 downto 0)  := (others => '0'); --                           .byteenable
		adapt_fir_mem_clk2_clk                     : in  std_logic                     := '0';             --         adapt_fir_mem_clk2.clk
		adapt_fir_mem_reset2_reset                 : in  std_logic                     := '0';             --       adapt_fir_mem_reset2.reset
		adapt_fir_mem_reset2_reset_req             : in  std_logic                     := '0';             --                           .reset_req
		micfilter_cntl_export                      : out std_logic_vector(31 downto 0);                    --             micfilter_cntl.export
		micfilter_rst_export                       : out std_logic;                                        --              micfilter_rst.export
		micfilter_adjust_export                    : out std_logic                                         --           micfilter_adjust.export
	);
end entity de2i_150_qsys;

architecture rtl of de2i_150_qsys is
	component de2i_150_qsys_pcie_ip is
		generic (
			p_pcie_hip_type                     : string                        := "0";
			lane_mask                           : std_logic_vector(7 downto 0)  := "00000000";
			max_link_width                      : integer                       := 4;
			millisecond_cycle_count             : string                        := "125000";
			enable_gen2_core                    : string                        := "false";
			gen2_lane_rate_mode                 : string                        := "false";
			no_soft_reset                       : string                        := "false";
			core_clk_divider                    : integer                       := 2;
			enable_ch0_pclk_out                 : string                        := "false";
			core_clk_source                     : string                        := "false";
			CB_P2A_AVALON_ADDR_B0               : integer                       := 0;
			bar0_size_mask                      : integer                       := 0;
			bar0_io_space                       : string                        := "false";
			bar0_64bit_mem_space                : string                        := "true";
			bar0_prefetchable                   : string                        := "true";
			CB_P2A_AVALON_ADDR_B1               : integer                       := 0;
			bar1_size_mask                      : integer                       := 0;
			bar1_io_space                       : string                        := "false";
			bar1_64bit_mem_space                : string                        := "true";
			bar1_prefetchable                   : string                        := "false";
			CB_P2A_AVALON_ADDR_B2               : integer                       := 0;
			bar2_size_mask                      : integer                       := 0;
			bar2_io_space                       : string                        := "false";
			bar2_64bit_mem_space                : string                        := "false";
			bar2_prefetchable                   : string                        := "false";
			CB_P2A_AVALON_ADDR_B3               : integer                       := 0;
			bar3_size_mask                      : integer                       := 0;
			bar3_io_space                       : string                        := "false";
			bar3_64bit_mem_space                : string                        := "false";
			bar3_prefetchable                   : string                        := "false";
			CB_P2A_AVALON_ADDR_B4               : integer                       := 0;
			bar4_size_mask                      : integer                       := 0;
			bar4_io_space                       : string                        := "false";
			bar4_64bit_mem_space                : string                        := "false";
			bar4_prefetchable                   : string                        := "false";
			CB_P2A_AVALON_ADDR_B5               : integer                       := 0;
			bar5_size_mask                      : integer                       := 0;
			bar5_io_space                       : string                        := "false";
			bar5_64bit_mem_space                : string                        := "false";
			bar5_prefetchable                   : string                        := "false";
			vendor_id                           : integer                       := 4466;
			device_id                           : integer                       := 4;
			revision_id                         : integer                       := 1;
			class_code                          : integer                       := 0;
			subsystem_vendor_id                 : integer                       := 4466;
			subsystem_device_id                 : integer                       := 4;
			port_link_number                    : integer                       := 1;
			msi_function_count                  : integer                       := 0;
			enable_msi_64bit_addressing         : string                        := "true";
			enable_function_msix_support        : string                        := "false";
			eie_before_nfts_count               : integer                       := 4;
			enable_completion_timeout_disable   : string                        := "false";
			completion_timeout                  : string                        := "NONE";
			enable_adapter_half_rate_mode       : string                        := "false";
			msix_pba_bir                        : integer                       := 0;
			msix_pba_offset                     : integer                       := 0;
			msix_table_bir                      : integer                       := 0;
			msix_table_offset                   : integer                       := 0;
			msix_table_size                     : integer                       := 0;
			use_crc_forwarding                  : string                        := "false";
			surprise_down_error_support         : string                        := "false";
			dll_active_report_support           : string                        := "false";
			bar_io_window_size                  : string                        := "32BIT";
			bar_prefetchable                    : integer                       := 32;
			hot_plug_support                    : std_logic_vector(6 downto 0)  := "0000000";
			no_command_completed                : string                        := "true";
			slot_power_limit                    : integer                       := 0;
			slot_power_scale                    : integer                       := 0;
			slot_number                         : integer                       := 0;
			enable_slot_register                : string                        := "false";
			advanced_errors                     : string                        := "false";
			enable_ecrc_check                   : string                        := "false";
			enable_ecrc_gen                     : string                        := "false";
			max_payload_size                    : integer                       := 0;
			retry_buffer_last_active_address    : integer                       := 2047;
			credit_buffer_allocation_aux        : string                        := "ABSOLUTE";
			vc0_rx_flow_ctrl_posted_header      : integer                       := 17;
			vc0_rx_flow_ctrl_posted_data        : integer                       := 91;
			vc0_rx_flow_ctrl_nonposted_header   : integer                       := 20;
			vc0_rx_flow_ctrl_nonposted_data     : integer                       := 0;
			vc0_rx_flow_ctrl_compl_header       : integer                       := 0;
			vc0_rx_flow_ctrl_compl_data         : integer                       := 0;
			RX_BUF                              : integer                       := 9;
			RH_NUM                              : integer                       := 7;
			G_TAG_NUM0                          : integer                       := 32;
			endpoint_l0_latency                 : integer                       := 0;
			endpoint_l1_latency                 : integer                       := 0;
			enable_l1_aspm                      : string                        := "false";
			l01_entry_latency                   : integer                       := 31;
			diffclock_nfts_count                : integer                       := 255;
			sameclock_nfts_count                : integer                       := 255;
			l1_exit_latency_sameclock           : integer                       := 7;
			l1_exit_latency_diffclock           : integer                       := 7;
			l0_exit_latency_sameclock           : integer                       := 7;
			l0_exit_latency_diffclock           : integer                       := 7;
			gen2_diffclock_nfts_count           : integer                       := 255;
			gen2_sameclock_nfts_count           : integer                       := 255;
			CG_COMMON_CLOCK_MODE                : integer                       := 1;
			CB_PCIE_MODE                        : integer                       := 0;
			AST_LITE                            : integer                       := 0;
			CB_PCIE_RX_LITE                     : integer                       := 0;
			CG_RXM_IRQ_NUM                      : integer                       := 16;
			CG_AVALON_S_ADDR_WIDTH              : integer                       := 20;
			bypass_tl                           : string                        := "false";
			CG_IMPL_CRA_AV_SLAVE_PORT           : integer                       := 1;
			CG_NO_CPL_REORDERING                : integer                       := 0;
			CG_ENABLE_A2P_INTERRUPT             : integer                       := 0;
			p_user_msi_enable                   : integer                       := 0;
			CG_IRQ_BIT_ENA                      : integer                       := 65535;
			CB_A2P_ADDR_MAP_IS_FIXED            : integer                       := 1;
			CB_A2P_ADDR_MAP_NUM_ENTRIES         : integer                       := 1;
			CB_A2P_ADDR_MAP_PASS_THRU_BITS      : integer                       := 20;
			CB_A2P_ADDR_MAP_FIXED_TABLE_0_HIGH  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_0_LOW   : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_1_HIGH  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_1_LOW   : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_2_HIGH  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_2_LOW   : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_3_HIGH  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_3_LOW   : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_4_HIGH  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_4_LOW   : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_5_HIGH  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_5_LOW   : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_6_HIGH  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_6_LOW   : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_7_HIGH  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_7_LOW   : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_8_HIGH  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_8_LOW   : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_9_HIGH  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_9_LOW   : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_10_HIGH : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_10_LOW  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_11_HIGH : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_11_LOW  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_12_HIGH : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_12_LOW  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_13_HIGH : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_13_LOW  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_14_HIGH : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_14_LOW  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_15_HIGH : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			CB_A2P_ADDR_MAP_FIXED_TABLE_15_LOW  : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
			RXM_DATA_WIDTH                      : integer                       := 64;
			RXM_BEN_WIDTH                       : integer                       := 8;
			TL_SELECTION                        : integer                       := 1;
			pcie_mode                           : string                        := "SHARED_MODE";
			single_rx_detect                    : integer                       := 4;
			enable_coreclk_out_half_rate        : string                        := "false";
			low_priority_vc                     : integer                       := 0;
			link_width                          : integer                       := 4;
			cyclone4                            : integer                       := 1
		);
		port (
			pcie_core_clk_clk                  : out std_logic;                                        -- clk
			pcie_core_reset_reset_n            : out std_logic;                                        -- reset_n
			cal_blk_clk_clk                    : in  std_logic                     := 'X';             -- clk
			txs_address                        : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			txs_chipselect                     : in  std_logic                     := 'X';             -- chipselect
			txs_byteenable                     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			txs_readdata                       : out std_logic_vector(63 downto 0);                    -- readdata
			txs_writedata                      : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			txs_read                           : in  std_logic                     := 'X';             -- read
			txs_write                          : in  std_logic                     := 'X';             -- write
			txs_burstcount                     : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- burstcount
			txs_readdatavalid                  : out std_logic;                                        -- readdatavalid
			txs_waitrequest                    : out std_logic;                                        -- waitrequest
			refclk_export                      : in  std_logic                     := 'X';             -- export
			test_in_test_in                    : in  std_logic_vector(39 downto 0) := (others => 'X'); -- test_in
			pcie_rstn_export                   : in  std_logic                     := 'X';             -- export
			clocks_sim_clk250_export           : out std_logic;                                        -- clk250_export
			clocks_sim_clk500_export           : out std_logic;                                        -- clk500_export
			clocks_sim_clk125_export           : out std_logic;                                        -- clk125_export
			reconfig_busy_busy_altgxb_reconfig : in  std_logic                     := 'X';             -- busy_altgxb_reconfig
			pipe_ext_pipe_mode                 : in  std_logic                     := 'X';             -- pipe_mode
			pipe_ext_phystatus_ext             : in  std_logic                     := 'X';             -- phystatus_ext
			pipe_ext_rate_ext                  : out std_logic;                                        -- rate_ext
			pipe_ext_powerdown_ext             : out std_logic_vector(1 downto 0);                     -- powerdown_ext
			pipe_ext_txdetectrx_ext            : out std_logic;                                        -- txdetectrx_ext
			pipe_ext_rxelecidle0_ext           : in  std_logic                     := 'X';             -- rxelecidle0_ext
			pipe_ext_rxdata0_ext               : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- rxdata0_ext
			pipe_ext_rxstatus0_ext             : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- rxstatus0_ext
			pipe_ext_rxvalid0_ext              : in  std_logic                     := 'X';             -- rxvalid0_ext
			pipe_ext_rxdatak0_ext              : in  std_logic                     := 'X';             -- rxdatak0_ext
			pipe_ext_txdata0_ext               : out std_logic_vector(7 downto 0);                     -- txdata0_ext
			pipe_ext_txdatak0_ext              : out std_logic;                                        -- txdatak0_ext
			pipe_ext_rxpolarity0_ext           : out std_logic;                                        -- rxpolarity0_ext
			pipe_ext_txcompl0_ext              : out std_logic;                                        -- txcompl0_ext
			pipe_ext_txelecidle0_ext           : out std_logic;                                        -- txelecidle0_ext
			powerdown_pll_powerdown            : in  std_logic                     := 'X';             -- pll_powerdown
			powerdown_gxb_powerdown            : in  std_logic                     := 'X';             -- gxb_powerdown
			bar1_0_address                     : out std_logic_vector(31 downto 0);                    -- address
			bar1_0_read                        : out std_logic;                                        -- read
			bar1_0_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			bar1_0_write                       : out std_logic;                                        -- write
			bar1_0_readdatavalid               : in  std_logic                     := 'X';             -- readdatavalid
			bar1_0_readdata                    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			bar1_0_writedata                   : out std_logic_vector(63 downto 0);                    -- writedata
			bar1_0_burstcount                  : out std_logic_vector(6 downto 0);                     -- burstcount
			bar1_0_byteenable                  : out std_logic_vector(7 downto 0);                     -- byteenable
			bar2_address                       : out std_logic_vector(31 downto 0);                    -- address
			bar2_read                          : out std_logic;                                        -- read
			bar2_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			bar2_write                         : out std_logic;                                        -- write
			bar2_readdatavalid                 : in  std_logic                     := 'X';             -- readdatavalid
			bar2_readdata                      : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			bar2_writedata                     : out std_logic_vector(63 downto 0);                    -- writedata
			bar2_burstcount                    : out std_logic_vector(6 downto 0);                     -- burstcount
			bar2_byteenable                    : out std_logic_vector(7 downto 0);                     -- byteenable
			cra_chipselect                     : in  std_logic                     := 'X';             -- chipselect
			cra_address                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			cra_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cra_read                           : in  std_logic                     := 'X';             -- read
			cra_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			cra_write                          : in  std_logic                     := 'X';             -- write
			cra_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cra_waitrequest                    : out std_logic;                                        -- waitrequest
			cra_irq_irq                        : out std_logic;                                        -- irq
			rxm_irq_irq                        : in  std_logic_vector(15 downto 0) := (others => 'X'); -- irq
			rx_in_rx_datain_0                  : in  std_logic                     := 'X';             -- rx_datain_0
			tx_out_tx_dataout_0                : out std_logic;                                        -- tx_dataout_0
			reconfig_togxb_data                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- data
			reconfig_gxbclk_clk                : in  std_logic                     := 'X';             -- clk
			reconfig_fromgxb_0_data            : out std_logic_vector(4 downto 0);                     -- data
			fixedclk_clk                       : in  std_logic                     := 'X'              -- clk
		);
	end component de2i_150_qsys_pcie_ip;

	component de2i_150_qsys_sgdma is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			m_read_readdata               : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			m_read_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			m_read_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			m_read_address                : out std_logic_vector(31 downto 0);                    -- address
			m_read_read                   : out std_logic;                                        -- read
			m_write_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			m_write_address               : out std_logic_vector(31 downto 0);                    -- address
			m_write_write                 : out std_logic;                                        -- write
			m_write_writedata             : out std_logic_vector(63 downto 0);                    -- writedata
			m_write_byteenable            : out std_logic_vector(7 downto 0)                      -- byteenable
		);
	end component de2i_150_qsys_sgdma;

	component de2i_150_qsys_fir_memory is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X'              -- reset_req
		);
	end component de2i_150_qsys_fir_memory;

	component de2i_150_qsys_led is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component de2i_150_qsys_led;

	component de2i_150_qsys_button is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component de2i_150_qsys_button;

	component de2i_150_qsys_fifo_memory is
		port (
			wrclock                          : in  std_logic                     := 'X';             -- clk
			reset_n                          : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata   : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write       : in  std_logic                     := 'X';             -- write
			avalonmm_write_slave_waitrequest : out std_logic;                                        -- waitrequest
			avalonmm_read_slave_readdata     : out std_logic_vector(63 downto 0);                    -- readdata
			avalonmm_read_slave_read         : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_waitrequest  : out std_logic;                                        -- waitrequest
			wrclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			wrclk_control_slave_irq          : out std_logic                                         -- irq
		);
	end component de2i_150_qsys_fifo_memory;

	component de2i_150_qsys_Interpo_4_0 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X'              -- reset_req
		);
	end component de2i_150_qsys_Interpo_4_0;

	component de2i_150_qsys_Interpo_5_0 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X'              -- reset_req
		);
	end component de2i_150_qsys_Interpo_5_0;

	component de2i_150_qsys_Interpo_5_1 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X'              -- reset_req
		);
	end component de2i_150_qsys_Interpo_5_1;

	component de2i_150_qsys_Interpo_5_2 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X'              -- reset_req
		);
	end component de2i_150_qsys_Interpo_5_2;

	component de2i_150_qsys_Interpo_5_3 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X'              -- reset_req
		);
	end component de2i_150_qsys_Interpo_5_3;

	component de2i_150_qsys_Adapt_FIR_mem is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X'              -- reset_req
		);
	end component de2i_150_qsys_Adapt_FIR_mem;

	component de2i_150_qsys_micFilter_cntl is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component de2i_150_qsys_micFilter_cntl;

	component de2i_150_qsys_micFilter_rst is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component de2i_150_qsys_micFilter_rst;

	component de2i_150_qsys_mm_interconnect_0 is
		port (
			pcie_ip_pcie_core_clk_clk                                   : in  std_logic                     := 'X';             -- clk
			pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			sgdma_reset_reset_bridge_in_reset_reset                     : in  std_logic                     := 'X';             -- reset
			pcie_ip_bar1_0_address                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			pcie_ip_bar1_0_waitrequest                                  : out std_logic;                                        -- waitrequest
			pcie_ip_bar1_0_burstcount                                   : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- burstcount
			pcie_ip_bar1_0_byteenable                                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			pcie_ip_bar1_0_read                                         : in  std_logic                     := 'X';             -- read
			pcie_ip_bar1_0_readdata                                     : out std_logic_vector(63 downto 0);                    -- readdata
			pcie_ip_bar1_0_readdatavalid                                : out std_logic;                                        -- readdatavalid
			pcie_ip_bar1_0_write                                        : in  std_logic                     := 'X';             -- write
			pcie_ip_bar1_0_writedata                                    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			sgdma_descriptor_read_address                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_descriptor_read_waitrequest                           : out std_logic;                                        -- waitrequest
			sgdma_descriptor_read_read                                  : in  std_logic                     := 'X';             -- read
			sgdma_descriptor_read_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_descriptor_read_readdatavalid                         : out std_logic;                                        -- readdatavalid
			sgdma_descriptor_write_address                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_descriptor_write_waitrequest                          : out std_logic;                                        -- waitrequest
			sgdma_descriptor_write_write                                : in  std_logic                     := 'X';             -- write
			sgdma_descriptor_write_writedata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_m_read_address                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_m_read_waitrequest                                    : out std_logic;                                        -- waitrequest
			sgdma_m_read_read                                           : in  std_logic                     := 'X';             -- read
			sgdma_m_read_readdata                                       : out std_logic_vector(63 downto 0);                    -- readdata
			sgdma_m_read_readdatavalid                                  : out std_logic;                                        -- readdatavalid
			sgdma_m_write_address                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_m_write_waitrequest                                   : out std_logic;                                        -- waitrequest
			sgdma_m_write_byteenable                                    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			sgdma_m_write_write                                         : in  std_logic                     := 'X';             -- write
			sgdma_m_write_writedata                                     : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			Adapt_FIR_mem_s1_address                                    : out std_logic_vector(8 downto 0);                     -- address
			Adapt_FIR_mem_s1_write                                      : out std_logic;                                        -- write
			Adapt_FIR_mem_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Adapt_FIR_mem_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			Adapt_FIR_mem_s1_byteenable                                 : out std_logic_vector(3 downto 0);                     -- byteenable
			Adapt_FIR_mem_s1_chipselect                                 : out std_logic;                                        -- chipselect
			Adapt_FIR_mem_s1_clken                                      : out std_logic;                                        -- clken
			button_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			button_s1_write                                             : out std_logic;                                        -- write
			button_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			button_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			button_s1_chipselect                                        : out std_logic;                                        -- chipselect
			fifo_memory_in_write                                        : out std_logic;                                        -- write
			fifo_memory_in_writedata                                    : out std_logic_vector(63 downto 0);                    -- writedata
			fifo_memory_in_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			fifo_memory_in_csr_address                                  : out std_logic_vector(2 downto 0);                     -- address
			fifo_memory_in_csr_write                                    : out std_logic;                                        -- write
			fifo_memory_in_csr_read                                     : out std_logic;                                        -- read
			fifo_memory_in_csr_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fifo_memory_in_csr_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			fifo_memory_out_read                                        : out std_logic;                                        -- read
			fifo_memory_out_readdata                                    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			fifo_memory_out_waitrequest                                 : in  std_logic                     := 'X';             -- waitrequest
			fir_memory_s1_address                                       : out std_logic_vector(9 downto 0);                     -- address
			fir_memory_s1_write                                         : out std_logic;                                        -- write
			fir_memory_s1_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			fir_memory_s1_writedata                                     : out std_logic_vector(31 downto 0);                    -- writedata
			fir_memory_s1_byteenable                                    : out std_logic_vector(3 downto 0);                     -- byteenable
			fir_memory_s1_chipselect                                    : out std_logic;                                        -- chipselect
			fir_memory_s1_clken                                         : out std_logic;                                        -- clken
			Interpo_4_0_s1_address                                      : out std_logic_vector(4 downto 0);                     -- address
			Interpo_4_0_s1_write                                        : out std_logic;                                        -- write
			Interpo_4_0_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Interpo_4_0_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			Interpo_4_0_s1_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			Interpo_4_0_s1_chipselect                                   : out std_logic;                                        -- chipselect
			Interpo_4_0_s1_clken                                        : out std_logic;                                        -- clken
			Interpo_5_0_s1_address                                      : out std_logic_vector(5 downto 0);                     -- address
			Interpo_5_0_s1_write                                        : out std_logic;                                        -- write
			Interpo_5_0_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Interpo_5_0_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			Interpo_5_0_s1_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			Interpo_5_0_s1_chipselect                                   : out std_logic;                                        -- chipselect
			Interpo_5_0_s1_clken                                        : out std_logic;                                        -- clken
			Interpo_5_1_s1_address                                      : out std_logic_vector(5 downto 0);                     -- address
			Interpo_5_1_s1_write                                        : out std_logic;                                        -- write
			Interpo_5_1_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Interpo_5_1_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			Interpo_5_1_s1_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			Interpo_5_1_s1_chipselect                                   : out std_logic;                                        -- chipselect
			Interpo_5_1_s1_clken                                        : out std_logic;                                        -- clken
			Interpo_5_2_s1_address                                      : out std_logic_vector(5 downto 0);                     -- address
			Interpo_5_2_s1_write                                        : out std_logic;                                        -- write
			Interpo_5_2_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Interpo_5_2_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			Interpo_5_2_s1_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			Interpo_5_2_s1_chipselect                                   : out std_logic;                                        -- chipselect
			Interpo_5_2_s1_clken                                        : out std_logic;                                        -- clken
			Interpo_5_3_s1_address                                      : out std_logic_vector(5 downto 0);                     -- address
			Interpo_5_3_s1_write                                        : out std_logic;                                        -- write
			Interpo_5_3_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Interpo_5_3_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			Interpo_5_3_s1_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			Interpo_5_3_s1_chipselect                                   : out std_logic;                                        -- chipselect
			Interpo_5_3_s1_clken                                        : out std_logic;                                        -- clken
			led_s1_address                                              : out std_logic_vector(1 downto 0);                     -- address
			led_s1_write                                                : out std_logic;                                        -- write
			led_s1_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_s1_writedata                                            : out std_logic_vector(31 downto 0);                    -- writedata
			led_s1_chipselect                                           : out std_logic;                                        -- chipselect
			micFilter_adjust_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			micFilter_adjust_s1_write                                   : out std_logic;                                        -- write
			micFilter_adjust_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			micFilter_adjust_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			micFilter_adjust_s1_chipselect                              : out std_logic;                                        -- chipselect
			micFilter_cntl_s1_address                                   : out std_logic_vector(2 downto 0);                     -- address
			micFilter_cntl_s1_write                                     : out std_logic;                                        -- write
			micFilter_cntl_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			micFilter_cntl_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			micFilter_cntl_s1_chipselect                                : out std_logic;                                        -- chipselect
			micFilter_rst_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			micFilter_rst_s1_write                                      : out std_logic;                                        -- write
			micFilter_rst_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			micFilter_rst_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			micFilter_rst_s1_chipselect                                 : out std_logic;                                        -- chipselect
			pcie_ip_txs_address                                         : out std_logic_vector(30 downto 0);                    -- address
			pcie_ip_txs_write                                           : out std_logic;                                        -- write
			pcie_ip_txs_read                                            : out std_logic;                                        -- read
			pcie_ip_txs_readdata                                        : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			pcie_ip_txs_writedata                                       : out std_logic_vector(63 downto 0);                    -- writedata
			pcie_ip_txs_burstcount                                      : out std_logic_vector(6 downto 0);                     -- burstcount
			pcie_ip_txs_byteenable                                      : out std_logic_vector(7 downto 0);                     -- byteenable
			pcie_ip_txs_readdatavalid                                   : in  std_logic                     := 'X';             -- readdatavalid
			pcie_ip_txs_waitrequest                                     : in  std_logic                     := 'X';             -- waitrequest
			pcie_ip_txs_chipselect                                      : out std_logic                                         -- chipselect
		);
	end component de2i_150_qsys_mm_interconnect_0;

	component de2i_150_qsys_mm_interconnect_1 is
		port (
			pcie_ip_pcie_core_clk_clk                                 : in  std_logic                     := 'X';             -- clk
			pcie_ip_bar2_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			sgdma_reset_reset_bridge_in_reset_reset                   : in  std_logic                     := 'X';             -- reset
			pcie_ip_bar2_address                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			pcie_ip_bar2_waitrequest                                  : out std_logic;                                        -- waitrequest
			pcie_ip_bar2_burstcount                                   : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- burstcount
			pcie_ip_bar2_byteenable                                   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			pcie_ip_bar2_read                                         : in  std_logic                     := 'X';             -- read
			pcie_ip_bar2_readdata                                     : out std_logic_vector(63 downto 0);                    -- readdata
			pcie_ip_bar2_readdatavalid                                : out std_logic;                                        -- readdatavalid
			pcie_ip_bar2_write                                        : in  std_logic                     := 'X';             -- write
			pcie_ip_bar2_writedata                                    : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			pcie_ip_cra_address                                       : out std_logic_vector(11 downto 0);                    -- address
			pcie_ip_cra_write                                         : out std_logic;                                        -- write
			pcie_ip_cra_read                                          : out std_logic;                                        -- read
			pcie_ip_cra_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pcie_ip_cra_writedata                                     : out std_logic_vector(31 downto 0);                    -- writedata
			pcie_ip_cra_byteenable                                    : out std_logic_vector(3 downto 0);                     -- byteenable
			pcie_ip_cra_waitrequest                                   : in  std_logic                     := 'X';             -- waitrequest
			pcie_ip_cra_chipselect                                    : out std_logic;                                        -- chipselect
			sgdma_csr_address                                         : out std_logic_vector(3 downto 0);                     -- address
			sgdma_csr_write                                           : out std_logic;                                        -- write
			sgdma_csr_read                                            : out std_logic;                                        -- read
			sgdma_csr_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_csr_writedata                                       : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_csr_chipselect                                      : out std_logic                                         -- chipselect
		);
	end component de2i_150_qsys_mm_interconnect_1;

	component de2i_150_qsys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(15 downto 0)         -- irq
		);
	end component de2i_150_qsys_irq_mapper;

	component de2i_150_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component de2i_150_qsys_rst_controller;

	component de2i_150_qsys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component de2i_150_qsys_rst_controller_001;

	signal pcie_ip_pcie_core_clk_clk                             : std_logic;                     -- pcie_ip:pcie_core_clk_clk -> [Adapt_FIR_mem:clk, Interpo_4_0:clk, Interpo_5_0:clk, Interpo_5_1:clk, Interpo_5_2:clk, Interpo_5_3:clk, button:clk, fifo_memory:wrclock, fir_memory:clk, irq_mapper:clk, led:clk, micFilter_adjust:clk, micFilter_cntl:clk, micFilter_rst:clk, mm_interconnect_0:pcie_ip_pcie_core_clk_clk, mm_interconnect_1:pcie_ip_pcie_core_clk_clk, pcie_ip:fixedclk_clk, rst_controller:clk, rst_controller_001:clk, sgdma:clk]
	signal pcie_ip_bar1_0_burstcount                             : std_logic_vector(6 downto 0);  -- pcie_ip:bar1_0_burstcount -> mm_interconnect_0:pcie_ip_bar1_0_burstcount
	signal pcie_ip_bar1_0_waitrequest                            : std_logic;                     -- mm_interconnect_0:pcie_ip_bar1_0_waitrequest -> pcie_ip:bar1_0_waitrequest
	signal pcie_ip_bar1_0_writedata                              : std_logic_vector(63 downto 0); -- pcie_ip:bar1_0_writedata -> mm_interconnect_0:pcie_ip_bar1_0_writedata
	signal pcie_ip_bar1_0_address                                : std_logic_vector(31 downto 0); -- pcie_ip:bar1_0_address -> mm_interconnect_0:pcie_ip_bar1_0_address
	signal pcie_ip_bar1_0_write                                  : std_logic;                     -- pcie_ip:bar1_0_write -> mm_interconnect_0:pcie_ip_bar1_0_write
	signal pcie_ip_bar1_0_read                                   : std_logic;                     -- pcie_ip:bar1_0_read -> mm_interconnect_0:pcie_ip_bar1_0_read
	signal pcie_ip_bar1_0_readdata                               : std_logic_vector(63 downto 0); -- mm_interconnect_0:pcie_ip_bar1_0_readdata -> pcie_ip:bar1_0_readdata
	signal pcie_ip_bar1_0_byteenable                             : std_logic_vector(7 downto 0);  -- pcie_ip:bar1_0_byteenable -> mm_interconnect_0:pcie_ip_bar1_0_byteenable
	signal pcie_ip_bar1_0_readdatavalid                          : std_logic;                     -- mm_interconnect_0:pcie_ip_bar1_0_readdatavalid -> pcie_ip:bar1_0_readdatavalid
	signal sgdma_m_read_waitrequest                              : std_logic;                     -- mm_interconnect_0:sgdma_m_read_waitrequest -> sgdma:m_read_waitrequest
	signal sgdma_m_read_address                                  : std_logic_vector(31 downto 0); -- sgdma:m_read_address -> mm_interconnect_0:sgdma_m_read_address
	signal sgdma_m_read_read                                     : std_logic;                     -- sgdma:m_read_read -> mm_interconnect_0:sgdma_m_read_read
	signal sgdma_m_read_readdata                                 : std_logic_vector(63 downto 0); -- mm_interconnect_0:sgdma_m_read_readdata -> sgdma:m_read_readdata
	signal sgdma_m_read_readdatavalid                            : std_logic;                     -- mm_interconnect_0:sgdma_m_read_readdatavalid -> sgdma:m_read_readdatavalid
	signal sgdma_m_write_waitrequest                             : std_logic;                     -- mm_interconnect_0:sgdma_m_write_waitrequest -> sgdma:m_write_waitrequest
	signal sgdma_m_write_writedata                               : std_logic_vector(63 downto 0); -- sgdma:m_write_writedata -> mm_interconnect_0:sgdma_m_write_writedata
	signal sgdma_m_write_address                                 : std_logic_vector(31 downto 0); -- sgdma:m_write_address -> mm_interconnect_0:sgdma_m_write_address
	signal sgdma_m_write_write                                   : std_logic;                     -- sgdma:m_write_write -> mm_interconnect_0:sgdma_m_write_write
	signal sgdma_m_write_byteenable                              : std_logic_vector(7 downto 0);  -- sgdma:m_write_byteenable -> mm_interconnect_0:sgdma_m_write_byteenable
	signal sgdma_descriptor_read_waitrequest                     : std_logic;                     -- mm_interconnect_0:sgdma_descriptor_read_waitrequest -> sgdma:descriptor_read_waitrequest
	signal sgdma_descriptor_read_address                         : std_logic_vector(31 downto 0); -- sgdma:descriptor_read_address -> mm_interconnect_0:sgdma_descriptor_read_address
	signal sgdma_descriptor_read_read                            : std_logic;                     -- sgdma:descriptor_read_read -> mm_interconnect_0:sgdma_descriptor_read_read
	signal sgdma_descriptor_read_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_descriptor_read_readdata -> sgdma:descriptor_read_readdata
	signal sgdma_descriptor_read_readdatavalid                   : std_logic;                     -- mm_interconnect_0:sgdma_descriptor_read_readdatavalid -> sgdma:descriptor_read_readdatavalid
	signal sgdma_descriptor_write_waitrequest                    : std_logic;                     -- mm_interconnect_0:sgdma_descriptor_write_waitrequest -> sgdma:descriptor_write_waitrequest
	signal sgdma_descriptor_write_writedata                      : std_logic_vector(31 downto 0); -- sgdma:descriptor_write_writedata -> mm_interconnect_0:sgdma_descriptor_write_writedata
	signal sgdma_descriptor_write_address                        : std_logic_vector(31 downto 0); -- sgdma:descriptor_write_address -> mm_interconnect_0:sgdma_descriptor_write_address
	signal sgdma_descriptor_write_write                          : std_logic;                     -- sgdma:descriptor_write_write -> mm_interconnect_0:sgdma_descriptor_write_write
	signal mm_interconnect_0_fir_memory_s1_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:fir_memory_s1_writedata -> fir_memory:writedata
	signal mm_interconnect_0_fir_memory_s1_address               : std_logic_vector(9 downto 0);  -- mm_interconnect_0:fir_memory_s1_address -> fir_memory:address
	signal mm_interconnect_0_fir_memory_s1_chipselect            : std_logic;                     -- mm_interconnect_0:fir_memory_s1_chipselect -> fir_memory:chipselect
	signal mm_interconnect_0_fir_memory_s1_clken                 : std_logic;                     -- mm_interconnect_0:fir_memory_s1_clken -> fir_memory:clken
	signal mm_interconnect_0_fir_memory_s1_write                 : std_logic;                     -- mm_interconnect_0:fir_memory_s1_write -> fir_memory:write
	signal mm_interconnect_0_fir_memory_s1_readdata              : std_logic_vector(31 downto 0); -- fir_memory:readdata -> mm_interconnect_0:fir_memory_s1_readdata
	signal mm_interconnect_0_fir_memory_s1_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:fir_memory_s1_byteenable -> fir_memory:byteenable
	signal mm_interconnect_0_led_s1_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_s1_writedata -> led:writedata
	signal mm_interconnect_0_led_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_s1_address -> led:address
	signal mm_interconnect_0_led_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:led_s1_chipselect -> led:chipselect
	signal mm_interconnect_0_led_s1_write                        : std_logic;                     -- mm_interconnect_0:led_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_readdata                     : std_logic_vector(31 downto 0); -- led:readdata -> mm_interconnect_0:led_s1_readdata
	signal mm_interconnect_0_button_s1_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:button_s1_writedata -> button:writedata
	signal mm_interconnect_0_button_s1_address                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button_s1_address -> button:address
	signal mm_interconnect_0_button_s1_chipselect                : std_logic;                     -- mm_interconnect_0:button_s1_chipselect -> button:chipselect
	signal mm_interconnect_0_button_s1_write                     : std_logic;                     -- mm_interconnect_0:button_s1_write -> mm_interconnect_0_button_s1_write:in
	signal mm_interconnect_0_button_s1_readdata                  : std_logic_vector(31 downto 0); -- button:readdata -> mm_interconnect_0:button_s1_readdata
	signal mm_interconnect_0_fifo_memory_in_csr_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:fifo_memory_in_csr_writedata -> fifo_memory:wrclk_control_slave_writedata
	signal mm_interconnect_0_fifo_memory_in_csr_address          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:fifo_memory_in_csr_address -> fifo_memory:wrclk_control_slave_address
	signal mm_interconnect_0_fifo_memory_in_csr_write            : std_logic;                     -- mm_interconnect_0:fifo_memory_in_csr_write -> fifo_memory:wrclk_control_slave_write
	signal mm_interconnect_0_fifo_memory_in_csr_read             : std_logic;                     -- mm_interconnect_0:fifo_memory_in_csr_read -> fifo_memory:wrclk_control_slave_read
	signal mm_interconnect_0_fifo_memory_in_csr_readdata         : std_logic_vector(31 downto 0); -- fifo_memory:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_memory_in_csr_readdata
	signal mm_interconnect_0_fifo_memory_in_waitrequest          : std_logic;                     -- fifo_memory:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_memory_in_waitrequest
	signal mm_interconnect_0_fifo_memory_in_writedata            : std_logic_vector(63 downto 0); -- mm_interconnect_0:fifo_memory_in_writedata -> fifo_memory:avalonmm_write_slave_writedata
	signal mm_interconnect_0_fifo_memory_in_write                : std_logic;                     -- mm_interconnect_0:fifo_memory_in_write -> fifo_memory:avalonmm_write_slave_write
	signal mm_interconnect_0_fifo_memory_out_waitrequest         : std_logic;                     -- fifo_memory:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_memory_out_waitrequest
	signal mm_interconnect_0_fifo_memory_out_read                : std_logic;                     -- mm_interconnect_0:fifo_memory_out_read -> fifo_memory:avalonmm_read_slave_read
	signal mm_interconnect_0_fifo_memory_out_readdata            : std_logic_vector(63 downto 0); -- fifo_memory:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_memory_out_readdata
	signal mm_interconnect_0_interpo_4_0_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:Interpo_4_0_s1_writedata -> Interpo_4_0:writedata
	signal mm_interconnect_0_interpo_4_0_s1_address              : std_logic_vector(4 downto 0);  -- mm_interconnect_0:Interpo_4_0_s1_address -> Interpo_4_0:address
	signal mm_interconnect_0_interpo_4_0_s1_chipselect           : std_logic;                     -- mm_interconnect_0:Interpo_4_0_s1_chipselect -> Interpo_4_0:chipselect
	signal mm_interconnect_0_interpo_4_0_s1_clken                : std_logic;                     -- mm_interconnect_0:Interpo_4_0_s1_clken -> Interpo_4_0:clken
	signal mm_interconnect_0_interpo_4_0_s1_write                : std_logic;                     -- mm_interconnect_0:Interpo_4_0_s1_write -> Interpo_4_0:write
	signal mm_interconnect_0_interpo_4_0_s1_readdata             : std_logic_vector(31 downto 0); -- Interpo_4_0:readdata -> mm_interconnect_0:Interpo_4_0_s1_readdata
	signal mm_interconnect_0_interpo_4_0_s1_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Interpo_4_0_s1_byteenable -> Interpo_4_0:byteenable
	signal mm_interconnect_0_interpo_5_0_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:Interpo_5_0_s1_writedata -> Interpo_5_0:writedata
	signal mm_interconnect_0_interpo_5_0_s1_address              : std_logic_vector(5 downto 0);  -- mm_interconnect_0:Interpo_5_0_s1_address -> Interpo_5_0:address
	signal mm_interconnect_0_interpo_5_0_s1_chipselect           : std_logic;                     -- mm_interconnect_0:Interpo_5_0_s1_chipselect -> Interpo_5_0:chipselect
	signal mm_interconnect_0_interpo_5_0_s1_clken                : std_logic;                     -- mm_interconnect_0:Interpo_5_0_s1_clken -> Interpo_5_0:clken
	signal mm_interconnect_0_interpo_5_0_s1_write                : std_logic;                     -- mm_interconnect_0:Interpo_5_0_s1_write -> Interpo_5_0:write
	signal mm_interconnect_0_interpo_5_0_s1_readdata             : std_logic_vector(31 downto 0); -- Interpo_5_0:readdata -> mm_interconnect_0:Interpo_5_0_s1_readdata
	signal mm_interconnect_0_interpo_5_0_s1_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Interpo_5_0_s1_byteenable -> Interpo_5_0:byteenable
	signal mm_interconnect_0_interpo_5_1_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:Interpo_5_1_s1_writedata -> Interpo_5_1:writedata
	signal mm_interconnect_0_interpo_5_1_s1_address              : std_logic_vector(5 downto 0);  -- mm_interconnect_0:Interpo_5_1_s1_address -> Interpo_5_1:address
	signal mm_interconnect_0_interpo_5_1_s1_chipselect           : std_logic;                     -- mm_interconnect_0:Interpo_5_1_s1_chipselect -> Interpo_5_1:chipselect
	signal mm_interconnect_0_interpo_5_1_s1_clken                : std_logic;                     -- mm_interconnect_0:Interpo_5_1_s1_clken -> Interpo_5_1:clken
	signal mm_interconnect_0_interpo_5_1_s1_write                : std_logic;                     -- mm_interconnect_0:Interpo_5_1_s1_write -> Interpo_5_1:write
	signal mm_interconnect_0_interpo_5_1_s1_readdata             : std_logic_vector(31 downto 0); -- Interpo_5_1:readdata -> mm_interconnect_0:Interpo_5_1_s1_readdata
	signal mm_interconnect_0_interpo_5_1_s1_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Interpo_5_1_s1_byteenable -> Interpo_5_1:byteenable
	signal mm_interconnect_0_interpo_5_2_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:Interpo_5_2_s1_writedata -> Interpo_5_2:writedata
	signal mm_interconnect_0_interpo_5_2_s1_address              : std_logic_vector(5 downto 0);  -- mm_interconnect_0:Interpo_5_2_s1_address -> Interpo_5_2:address
	signal mm_interconnect_0_interpo_5_2_s1_chipselect           : std_logic;                     -- mm_interconnect_0:Interpo_5_2_s1_chipselect -> Interpo_5_2:chipselect
	signal mm_interconnect_0_interpo_5_2_s1_clken                : std_logic;                     -- mm_interconnect_0:Interpo_5_2_s1_clken -> Interpo_5_2:clken
	signal mm_interconnect_0_interpo_5_2_s1_write                : std_logic;                     -- mm_interconnect_0:Interpo_5_2_s1_write -> Interpo_5_2:write
	signal mm_interconnect_0_interpo_5_2_s1_readdata             : std_logic_vector(31 downto 0); -- Interpo_5_2:readdata -> mm_interconnect_0:Interpo_5_2_s1_readdata
	signal mm_interconnect_0_interpo_5_2_s1_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Interpo_5_2_s1_byteenable -> Interpo_5_2:byteenable
	signal mm_interconnect_0_interpo_5_3_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:Interpo_5_3_s1_writedata -> Interpo_5_3:writedata
	signal mm_interconnect_0_interpo_5_3_s1_address              : std_logic_vector(5 downto 0);  -- mm_interconnect_0:Interpo_5_3_s1_address -> Interpo_5_3:address
	signal mm_interconnect_0_interpo_5_3_s1_chipselect           : std_logic;                     -- mm_interconnect_0:Interpo_5_3_s1_chipselect -> Interpo_5_3:chipselect
	signal mm_interconnect_0_interpo_5_3_s1_clken                : std_logic;                     -- mm_interconnect_0:Interpo_5_3_s1_clken -> Interpo_5_3:clken
	signal mm_interconnect_0_interpo_5_3_s1_write                : std_logic;                     -- mm_interconnect_0:Interpo_5_3_s1_write -> Interpo_5_3:write
	signal mm_interconnect_0_interpo_5_3_s1_readdata             : std_logic_vector(31 downto 0); -- Interpo_5_3:readdata -> mm_interconnect_0:Interpo_5_3_s1_readdata
	signal mm_interconnect_0_interpo_5_3_s1_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Interpo_5_3_s1_byteenable -> Interpo_5_3:byteenable
	signal mm_interconnect_0_adapt_fir_mem_s1_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:Adapt_FIR_mem_s1_writedata -> Adapt_FIR_mem:writedata
	signal mm_interconnect_0_adapt_fir_mem_s1_address            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:Adapt_FIR_mem_s1_address -> Adapt_FIR_mem:address
	signal mm_interconnect_0_adapt_fir_mem_s1_chipselect         : std_logic;                     -- mm_interconnect_0:Adapt_FIR_mem_s1_chipselect -> Adapt_FIR_mem:chipselect
	signal mm_interconnect_0_adapt_fir_mem_s1_clken              : std_logic;                     -- mm_interconnect_0:Adapt_FIR_mem_s1_clken -> Adapt_FIR_mem:clken
	signal mm_interconnect_0_adapt_fir_mem_s1_write              : std_logic;                     -- mm_interconnect_0:Adapt_FIR_mem_s1_write -> Adapt_FIR_mem:write
	signal mm_interconnect_0_adapt_fir_mem_s1_readdata           : std_logic_vector(31 downto 0); -- Adapt_FIR_mem:readdata -> mm_interconnect_0:Adapt_FIR_mem_s1_readdata
	signal mm_interconnect_0_adapt_fir_mem_s1_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Adapt_FIR_mem_s1_byteenable -> Adapt_FIR_mem:byteenable
	signal mm_interconnect_0_micfilter_cntl_s1_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:micFilter_cntl_s1_writedata -> micFilter_cntl:writedata
	signal mm_interconnect_0_micfilter_cntl_s1_address           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:micFilter_cntl_s1_address -> micFilter_cntl:address
	signal mm_interconnect_0_micfilter_cntl_s1_chipselect        : std_logic;                     -- mm_interconnect_0:micFilter_cntl_s1_chipselect -> micFilter_cntl:chipselect
	signal mm_interconnect_0_micfilter_cntl_s1_write             : std_logic;                     -- mm_interconnect_0:micFilter_cntl_s1_write -> mm_interconnect_0_micfilter_cntl_s1_write:in
	signal mm_interconnect_0_micfilter_cntl_s1_readdata          : std_logic_vector(31 downto 0); -- micFilter_cntl:readdata -> mm_interconnect_0:micFilter_cntl_s1_readdata
	signal mm_interconnect_0_micfilter_rst_s1_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:micFilter_rst_s1_writedata -> micFilter_rst:writedata
	signal mm_interconnect_0_micfilter_rst_s1_address            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:micFilter_rst_s1_address -> micFilter_rst:address
	signal mm_interconnect_0_micfilter_rst_s1_chipselect         : std_logic;                     -- mm_interconnect_0:micFilter_rst_s1_chipselect -> micFilter_rst:chipselect
	signal mm_interconnect_0_micfilter_rst_s1_write              : std_logic;                     -- mm_interconnect_0:micFilter_rst_s1_write -> mm_interconnect_0_micfilter_rst_s1_write:in
	signal mm_interconnect_0_micfilter_rst_s1_readdata           : std_logic_vector(31 downto 0); -- micFilter_rst:readdata -> mm_interconnect_0:micFilter_rst_s1_readdata
	signal mm_interconnect_0_micfilter_adjust_s1_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:micFilter_adjust_s1_writedata -> micFilter_adjust:writedata
	signal mm_interconnect_0_micfilter_adjust_s1_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:micFilter_adjust_s1_address -> micFilter_adjust:address
	signal mm_interconnect_0_micfilter_adjust_s1_chipselect      : std_logic;                     -- mm_interconnect_0:micFilter_adjust_s1_chipselect -> micFilter_adjust:chipselect
	signal mm_interconnect_0_micfilter_adjust_s1_write           : std_logic;                     -- mm_interconnect_0:micFilter_adjust_s1_write -> mm_interconnect_0_micfilter_adjust_s1_write:in
	signal mm_interconnect_0_micfilter_adjust_s1_readdata        : std_logic_vector(31 downto 0); -- micFilter_adjust:readdata -> mm_interconnect_0:micFilter_adjust_s1_readdata
	signal mm_interconnect_0_pcie_ip_txs_waitrequest             : std_logic;                     -- pcie_ip:txs_waitrequest -> mm_interconnect_0:pcie_ip_txs_waitrequest
	signal mm_interconnect_0_pcie_ip_txs_burstcount              : std_logic_vector(6 downto 0);  -- mm_interconnect_0:pcie_ip_txs_burstcount -> pcie_ip:txs_burstcount
	signal mm_interconnect_0_pcie_ip_txs_writedata               : std_logic_vector(63 downto 0); -- mm_interconnect_0:pcie_ip_txs_writedata -> pcie_ip:txs_writedata
	signal mm_interconnect_0_pcie_ip_txs_address                 : std_logic_vector(30 downto 0); -- mm_interconnect_0:pcie_ip_txs_address -> pcie_ip:txs_address
	signal mm_interconnect_0_pcie_ip_txs_chipselect              : std_logic;                     -- mm_interconnect_0:pcie_ip_txs_chipselect -> pcie_ip:txs_chipselect
	signal mm_interconnect_0_pcie_ip_txs_write                   : std_logic;                     -- mm_interconnect_0:pcie_ip_txs_write -> pcie_ip:txs_write
	signal mm_interconnect_0_pcie_ip_txs_read                    : std_logic;                     -- mm_interconnect_0:pcie_ip_txs_read -> pcie_ip:txs_read
	signal mm_interconnect_0_pcie_ip_txs_readdata                : std_logic_vector(63 downto 0); -- pcie_ip:txs_readdata -> mm_interconnect_0:pcie_ip_txs_readdata
	signal mm_interconnect_0_pcie_ip_txs_readdatavalid           : std_logic;                     -- pcie_ip:txs_readdatavalid -> mm_interconnect_0:pcie_ip_txs_readdatavalid
	signal mm_interconnect_0_pcie_ip_txs_byteenable              : std_logic_vector(7 downto 0);  -- mm_interconnect_0:pcie_ip_txs_byteenable -> pcie_ip:txs_byteenable
	signal pcie_ip_bar2_burstcount                               : std_logic_vector(6 downto 0);  -- pcie_ip:bar2_burstcount -> mm_interconnect_1:pcie_ip_bar2_burstcount
	signal pcie_ip_bar2_waitrequest                              : std_logic;                     -- mm_interconnect_1:pcie_ip_bar2_waitrequest -> pcie_ip:bar2_waitrequest
	signal pcie_ip_bar2_writedata                                : std_logic_vector(63 downto 0); -- pcie_ip:bar2_writedata -> mm_interconnect_1:pcie_ip_bar2_writedata
	signal pcie_ip_bar2_address                                  : std_logic_vector(31 downto 0); -- pcie_ip:bar2_address -> mm_interconnect_1:pcie_ip_bar2_address
	signal pcie_ip_bar2_write                                    : std_logic;                     -- pcie_ip:bar2_write -> mm_interconnect_1:pcie_ip_bar2_write
	signal pcie_ip_bar2_read                                     : std_logic;                     -- pcie_ip:bar2_read -> mm_interconnect_1:pcie_ip_bar2_read
	signal pcie_ip_bar2_readdata                                 : std_logic_vector(63 downto 0); -- mm_interconnect_1:pcie_ip_bar2_readdata -> pcie_ip:bar2_readdata
	signal pcie_ip_bar2_byteenable                               : std_logic_vector(7 downto 0);  -- pcie_ip:bar2_byteenable -> mm_interconnect_1:pcie_ip_bar2_byteenable
	signal pcie_ip_bar2_readdatavalid                            : std_logic;                     -- mm_interconnect_1:pcie_ip_bar2_readdatavalid -> pcie_ip:bar2_readdatavalid
	signal mm_interconnect_1_sgdma_csr_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_1:sgdma_csr_writedata -> sgdma:csr_writedata
	signal mm_interconnect_1_sgdma_csr_address                   : std_logic_vector(3 downto 0);  -- mm_interconnect_1:sgdma_csr_address -> sgdma:csr_address
	signal mm_interconnect_1_sgdma_csr_chipselect                : std_logic;                     -- mm_interconnect_1:sgdma_csr_chipselect -> sgdma:csr_chipselect
	signal mm_interconnect_1_sgdma_csr_write                     : std_logic;                     -- mm_interconnect_1:sgdma_csr_write -> sgdma:csr_write
	signal mm_interconnect_1_sgdma_csr_read                      : std_logic;                     -- mm_interconnect_1:sgdma_csr_read -> sgdma:csr_read
	signal mm_interconnect_1_sgdma_csr_readdata                  : std_logic_vector(31 downto 0); -- sgdma:csr_readdata -> mm_interconnect_1:sgdma_csr_readdata
	signal mm_interconnect_1_pcie_ip_cra_waitrequest             : std_logic;                     -- pcie_ip:cra_waitrequest -> mm_interconnect_1:pcie_ip_cra_waitrequest
	signal mm_interconnect_1_pcie_ip_cra_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_1:pcie_ip_cra_writedata -> pcie_ip:cra_writedata
	signal mm_interconnect_1_pcie_ip_cra_address                 : std_logic_vector(11 downto 0); -- mm_interconnect_1:pcie_ip_cra_address -> pcie_ip:cra_address
	signal mm_interconnect_1_pcie_ip_cra_chipselect              : std_logic;                     -- mm_interconnect_1:pcie_ip_cra_chipselect -> pcie_ip:cra_chipselect
	signal mm_interconnect_1_pcie_ip_cra_write                   : std_logic;                     -- mm_interconnect_1:pcie_ip_cra_write -> pcie_ip:cra_write
	signal mm_interconnect_1_pcie_ip_cra_read                    : std_logic;                     -- mm_interconnect_1:pcie_ip_cra_read -> pcie_ip:cra_read
	signal mm_interconnect_1_pcie_ip_cra_readdata                : std_logic_vector(31 downto 0); -- pcie_ip:cra_readdata -> mm_interconnect_1:pcie_ip_cra_readdata
	signal mm_interconnect_1_pcie_ip_cra_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_1:pcie_ip_cra_byteenable -> pcie_ip:cra_byteenable
	signal irq_mapper_receiver0_irq                              : std_logic;                     -- sgdma:csr_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                              : std_logic;                     -- fifo_memory:wrclk_control_slave_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                              : std_logic;                     -- button:irq -> irq_mapper:receiver2_irq
	signal pcie_ip_rxm_irq_irq                                   : std_logic_vector(15 downto 0); -- irq_mapper:sender_irq -> pcie_ip:rxm_irq_irq
	signal rst_controller_reset_out_reset                        : std_logic;                     -- rst_controller:reset_out -> [Adapt_FIR_mem:reset, Interpo_4_0:reset, Interpo_5_0:reset, Interpo_5_1:reset, Interpo_5_2:reset, Interpo_5_3:reset, fir_memory:reset, mm_interconnect_0:sgdma_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sgdma_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                    : std_logic;                     -- rst_controller:reset_req -> [Adapt_FIR_mem:reset_req, Interpo_4_0:reset_req, Interpo_5_0:reset_req, Interpo_5_1:reset_req, Interpo_5_2:reset_req, Interpo_5_3:reset_req, fir_memory:reset_req, rst_translator:reset_req_in]
	signal pcie_ip_pcie_core_reset_reset                         : std_logic;                     -- pcie_ip:pcie_core_reset_reset_n -> pcie_ip_pcie_core_reset_reset:in
	signal rst_controller_001_reset_out_reset                    : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pcie_ip_bar2_translator_reset_reset_bridge_in_reset_reset]
	signal reset_reset_n_ports_inv                               : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in1
	signal mm_interconnect_0_led_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> led:write_n
	signal mm_interconnect_0_button_s1_write_ports_inv           : std_logic;                     -- mm_interconnect_0_button_s1_write:inv -> button:write_n
	signal mm_interconnect_0_micfilter_cntl_s1_write_ports_inv   : std_logic;                     -- mm_interconnect_0_micfilter_cntl_s1_write:inv -> micFilter_cntl:write_n
	signal mm_interconnect_0_micfilter_rst_s1_write_ports_inv    : std_logic;                     -- mm_interconnect_0_micfilter_rst_s1_write:inv -> micFilter_rst:write_n
	signal mm_interconnect_0_micfilter_adjust_s1_write_ports_inv : std_logic;                     -- mm_interconnect_0_micfilter_adjust_s1_write:inv -> micFilter_adjust:write_n
	signal rst_controller_reset_out_reset_ports_inv              : std_logic;                     -- rst_controller_reset_out_reset:inv -> [button:reset_n, fifo_memory:reset_n, led:reset_n, micFilter_adjust:reset_n, micFilter_cntl:reset_n, micFilter_rst:reset_n, sgdma:system_reset_n]
	signal pcie_ip_pcie_core_reset_reset_ports_inv               : std_logic;                     -- pcie_ip_pcie_core_reset_reset:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]

begin

	pcie_ip : component de2i_150_qsys_pcie_ip
		generic map (
			p_pcie_hip_type                     => "2",
			lane_mask                           => "11111110",
			max_link_width                      => 1,
			millisecond_cycle_count             => "125000",
			enable_gen2_core                    => "false",
			gen2_lane_rate_mode                 => "false",
			no_soft_reset                       => "false",
			core_clk_divider                    => 2,
			enable_ch0_pclk_out                 => "true",
			core_clk_source                     => "pclk",
			CB_P2A_AVALON_ADDR_B0               => 0,
			bar0_size_mask                      => 19,
			bar0_io_space                       => "false",
			bar0_64bit_mem_space                => "true",
			bar0_prefetchable                   => "true",
			CB_P2A_AVALON_ADDR_B1               => 0,
			bar1_size_mask                      => 0,
			bar1_io_space                       => "false",
			bar1_64bit_mem_space                => "true",
			bar1_prefetchable                   => "false",
			CB_P2A_AVALON_ADDR_B2               => 0,
			bar2_size_mask                      => 15,
			bar2_io_space                       => "false",
			bar2_64bit_mem_space                => "false",
			bar2_prefetchable                   => "false",
			CB_P2A_AVALON_ADDR_B3               => 0,
			bar3_size_mask                      => 0,
			bar3_io_space                       => "false",
			bar3_64bit_mem_space                => "false",
			bar3_prefetchable                   => "false",
			CB_P2A_AVALON_ADDR_B4               => 0,
			bar4_size_mask                      => 0,
			bar4_io_space                       => "false",
			bar4_64bit_mem_space                => "false",
			bar4_prefetchable                   => "false",
			CB_P2A_AVALON_ADDR_B5               => 0,
			bar5_size_mask                      => 0,
			bar5_io_space                       => "false",
			bar5_64bit_mem_space                => "false",
			bar5_prefetchable                   => "false",
			vendor_id                           => 4466,
			device_id                           => 57345,
			revision_id                         => 1,
			class_code                          => 0,
			subsystem_vendor_id                 => 4466,
			subsystem_device_id                 => 4,
			port_link_number                    => 1,
			msi_function_count                  => 0,
			enable_msi_64bit_addressing         => "true",
			enable_function_msix_support        => "false",
			eie_before_nfts_count               => 4,
			enable_completion_timeout_disable   => "false",
			completion_timeout                  => "NONE",
			enable_adapter_half_rate_mode       => "false",
			msix_pba_bir                        => 0,
			msix_pba_offset                     => 0,
			msix_table_bir                      => 0,
			msix_table_offset                   => 0,
			msix_table_size                     => 0,
			use_crc_forwarding                  => "false",
			surprise_down_error_support         => "false",
			dll_active_report_support           => "false",
			bar_io_window_size                  => "32BIT",
			bar_prefetchable                    => 32,
			hot_plug_support                    => "0000000",
			no_command_completed                => "true",
			slot_power_limit                    => 0,
			slot_power_scale                    => 0,
			slot_number                         => 0,
			enable_slot_register                => "false",
			advanced_errors                     => "false",
			enable_ecrc_check                   => "false",
			enable_ecrc_gen                     => "false",
			max_payload_size                    => 0,
			retry_buffer_last_active_address    => 255,
			credit_buffer_allocation_aux        => "ABSOLUTE",
			vc0_rx_flow_ctrl_posted_header      => 28,
			vc0_rx_flow_ctrl_posted_data        => 198,
			vc0_rx_flow_ctrl_nonposted_header   => 30,
			vc0_rx_flow_ctrl_nonposted_data     => 0,
			vc0_rx_flow_ctrl_compl_header       => 48,
			vc0_rx_flow_ctrl_compl_data         => 256,
			RX_BUF                              => 9,
			RH_NUM                              => 7,
			G_TAG_NUM0                          => 32,
			endpoint_l0_latency                 => 0,
			endpoint_l1_latency                 => 0,
			enable_l1_aspm                      => "false",
			l01_entry_latency                   => 31,
			diffclock_nfts_count                => 255,
			sameclock_nfts_count                => 255,
			l1_exit_latency_sameclock           => 7,
			l1_exit_latency_diffclock           => 7,
			l0_exit_latency_sameclock           => 7,
			l0_exit_latency_diffclock           => 7,
			gen2_diffclock_nfts_count           => 255,
			gen2_sameclock_nfts_count           => 255,
			CG_COMMON_CLOCK_MODE                => 1,
			CB_PCIE_MODE                        => 0,
			AST_LITE                            => 0,
			CB_PCIE_RX_LITE                     => 0,
			CG_RXM_IRQ_NUM                      => 16,
			CG_AVALON_S_ADDR_WIDTH              => 20,
			bypass_tl                           => "false",
			CG_IMPL_CRA_AV_SLAVE_PORT           => 1,
			CG_NO_CPL_REORDERING                => 0,
			CG_ENABLE_A2P_INTERRUPT             => 0,
			p_user_msi_enable                   => 0,
			CG_IRQ_BIT_ENA                      => 65535,
			CB_A2P_ADDR_MAP_IS_FIXED            => 1,
			CB_A2P_ADDR_MAP_NUM_ENTRIES         => 1,
			CB_A2P_ADDR_MAP_PASS_THRU_BITS      => 31,
			CB_A2P_ADDR_MAP_FIXED_TABLE_0_HIGH  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_0_LOW   => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_1_HIGH  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_1_LOW   => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_2_HIGH  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_2_LOW   => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_3_HIGH  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_3_LOW   => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_4_HIGH  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_4_LOW   => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_5_HIGH  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_5_LOW   => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_6_HIGH  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_6_LOW   => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_7_HIGH  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_7_LOW   => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_8_HIGH  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_8_LOW   => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_9_HIGH  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_9_LOW   => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_10_HIGH => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_10_LOW  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_11_HIGH => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_11_LOW  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_12_HIGH => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_12_LOW  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_13_HIGH => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_13_LOW  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_14_HIGH => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_14_LOW  => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_15_HIGH => "00000000000000000000000000000000",
			CB_A2P_ADDR_MAP_FIXED_TABLE_15_LOW  => "00000000000000000000000000000000",
			RXM_DATA_WIDTH                      => 64,
			RXM_BEN_WIDTH                       => 8,
			TL_SELECTION                        => 1,
			pcie_mode                           => "SHARED_MODE",
			single_rx_detect                    => 1,
			enable_coreclk_out_half_rate        => "false",
			low_priority_vc                     => 0,
			link_width                          => 1,
			cyclone4                            => 1
		)
		port map (
			pcie_core_clk_clk                  => pcie_ip_pcie_core_clk_clk,                   --      pcie_core_clk.clk
			pcie_core_reset_reset_n            => pcie_ip_pcie_core_reset_reset,               --    pcie_core_reset.reset_n
			cal_blk_clk_clk                    => clk_clk,                                     --        cal_blk_clk.clk
			txs_address                        => mm_interconnect_0_pcie_ip_txs_address,       --                txs.address
			txs_chipselect                     => mm_interconnect_0_pcie_ip_txs_chipselect,    --                   .chipselect
			txs_byteenable                     => mm_interconnect_0_pcie_ip_txs_byteenable,    --                   .byteenable
			txs_readdata                       => mm_interconnect_0_pcie_ip_txs_readdata,      --                   .readdata
			txs_writedata                      => mm_interconnect_0_pcie_ip_txs_writedata,     --                   .writedata
			txs_read                           => mm_interconnect_0_pcie_ip_txs_read,          --                   .read
			txs_write                          => mm_interconnect_0_pcie_ip_txs_write,         --                   .write
			txs_burstcount                     => mm_interconnect_0_pcie_ip_txs_burstcount,    --                   .burstcount
			txs_readdatavalid                  => mm_interconnect_0_pcie_ip_txs_readdatavalid, --                   .readdatavalid
			txs_waitrequest                    => mm_interconnect_0_pcie_ip_txs_waitrequest,   --                   .waitrequest
			refclk_export                      => pcie_ip_refclk_export,                       --             refclk.export
			test_in_test_in                    => pcie_ip_test_in_test_in,                     --            test_in.test_in
			pcie_rstn_export                   => pcie_ip_pcie_rstn_export,                    --          pcie_rstn.export
			clocks_sim_clk250_export           => pcie_ip_clocks_sim_clk250_export,            --         clocks_sim.clk250_export
			clocks_sim_clk500_export           => pcie_ip_clocks_sim_clk500_export,            --                   .clk500_export
			clocks_sim_clk125_export           => pcie_ip_clocks_sim_clk125_export,            --                   .clk125_export
			reconfig_busy_busy_altgxb_reconfig => pcie_ip_reconfig_busy_busy_altgxb_reconfig,  --      reconfig_busy.busy_altgxb_reconfig
			pipe_ext_pipe_mode                 => pcie_ip_pipe_ext_pipe_mode,                  --           pipe_ext.pipe_mode
			pipe_ext_phystatus_ext             => pcie_ip_pipe_ext_phystatus_ext,              --                   .phystatus_ext
			pipe_ext_rate_ext                  => pcie_ip_pipe_ext_rate_ext,                   --                   .rate_ext
			pipe_ext_powerdown_ext             => pcie_ip_pipe_ext_powerdown_ext,              --                   .powerdown_ext
			pipe_ext_txdetectrx_ext            => pcie_ip_pipe_ext_txdetectrx_ext,             --                   .txdetectrx_ext
			pipe_ext_rxelecidle0_ext           => pcie_ip_pipe_ext_rxelecidle0_ext,            --                   .rxelecidle0_ext
			pipe_ext_rxdata0_ext               => pcie_ip_pipe_ext_rxdata0_ext,                --                   .rxdata0_ext
			pipe_ext_rxstatus0_ext             => pcie_ip_pipe_ext_rxstatus0_ext,              --                   .rxstatus0_ext
			pipe_ext_rxvalid0_ext              => pcie_ip_pipe_ext_rxvalid0_ext,               --                   .rxvalid0_ext
			pipe_ext_rxdatak0_ext              => pcie_ip_pipe_ext_rxdatak0_ext,               --                   .rxdatak0_ext
			pipe_ext_txdata0_ext               => pcie_ip_pipe_ext_txdata0_ext,                --                   .txdata0_ext
			pipe_ext_txdatak0_ext              => pcie_ip_pipe_ext_txdatak0_ext,               --                   .txdatak0_ext
			pipe_ext_rxpolarity0_ext           => pcie_ip_pipe_ext_rxpolarity0_ext,            --                   .rxpolarity0_ext
			pipe_ext_txcompl0_ext              => pcie_ip_pipe_ext_txcompl0_ext,               --                   .txcompl0_ext
			pipe_ext_txelecidle0_ext           => pcie_ip_pipe_ext_txelecidle0_ext,            --                   .txelecidle0_ext
			powerdown_pll_powerdown            => open,                                        --          powerdown.pll_powerdown
			powerdown_gxb_powerdown            => open,                                        --                   .gxb_powerdown
			bar1_0_address                     => pcie_ip_bar1_0_address,                      --             bar1_0.address
			bar1_0_read                        => pcie_ip_bar1_0_read,                         --                   .read
			bar1_0_waitrequest                 => pcie_ip_bar1_0_waitrequest,                  --                   .waitrequest
			bar1_0_write                       => pcie_ip_bar1_0_write,                        --                   .write
			bar1_0_readdatavalid               => pcie_ip_bar1_0_readdatavalid,                --                   .readdatavalid
			bar1_0_readdata                    => pcie_ip_bar1_0_readdata,                     --                   .readdata
			bar1_0_writedata                   => pcie_ip_bar1_0_writedata,                    --                   .writedata
			bar1_0_burstcount                  => pcie_ip_bar1_0_burstcount,                   --                   .burstcount
			bar1_0_byteenable                  => pcie_ip_bar1_0_byteenable,                   --                   .byteenable
			bar2_address                       => pcie_ip_bar2_address,                        --               bar2.address
			bar2_read                          => pcie_ip_bar2_read,                           --                   .read
			bar2_waitrequest                   => pcie_ip_bar2_waitrequest,                    --                   .waitrequest
			bar2_write                         => pcie_ip_bar2_write,                          --                   .write
			bar2_readdatavalid                 => pcie_ip_bar2_readdatavalid,                  --                   .readdatavalid
			bar2_readdata                      => pcie_ip_bar2_readdata,                       --                   .readdata
			bar2_writedata                     => pcie_ip_bar2_writedata,                      --                   .writedata
			bar2_burstcount                    => pcie_ip_bar2_burstcount,                     --                   .burstcount
			bar2_byteenable                    => pcie_ip_bar2_byteenable,                     --                   .byteenable
			cra_chipselect                     => mm_interconnect_1_pcie_ip_cra_chipselect,    --                cra.chipselect
			cra_address                        => mm_interconnect_1_pcie_ip_cra_address,       --                   .address
			cra_byteenable                     => mm_interconnect_1_pcie_ip_cra_byteenable,    --                   .byteenable
			cra_read                           => mm_interconnect_1_pcie_ip_cra_read,          --                   .read
			cra_readdata                       => mm_interconnect_1_pcie_ip_cra_readdata,      --                   .readdata
			cra_write                          => mm_interconnect_1_pcie_ip_cra_write,         --                   .write
			cra_writedata                      => mm_interconnect_1_pcie_ip_cra_writedata,     --                   .writedata
			cra_waitrequest                    => mm_interconnect_1_pcie_ip_cra_waitrequest,   --                   .waitrequest
			cra_irq_irq                        => open,                                        --            cra_irq.irq
			rxm_irq_irq                        => pcie_ip_rxm_irq_irq,                         --            rxm_irq.irq
			rx_in_rx_datain_0                  => pcie_ip_rx_in_rx_datain_0,                   --              rx_in.rx_datain_0
			tx_out_tx_dataout_0                => pcie_ip_tx_out_tx_dataout_0,                 --             tx_out.tx_dataout_0
			reconfig_togxb_data                => pcie_ip_reconfig_togxb_data,                 --     reconfig_togxb.data
			reconfig_gxbclk_clk                => clk_clk,                                     --    reconfig_gxbclk.clk
			reconfig_fromgxb_0_data            => pcie_ip_reconfig_fromgxb_0_data,             -- reconfig_fromgxb_0.data
			fixedclk_clk                       => pcie_ip_pcie_core_clk_clk                    --           fixedclk.clk
		);

	sgdma : component de2i_150_qsys_sgdma
		port map (
			clk                           => pcie_ip_pcie_core_clk_clk,                --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv, --            reset.reset_n
			csr_chipselect                => mm_interconnect_1_sgdma_csr_chipselect,   --              csr.chipselect
			csr_address                   => mm_interconnect_1_sgdma_csr_address,      --                 .address
			csr_read                      => mm_interconnect_1_sgdma_csr_read,         --                 .read
			csr_write                     => mm_interconnect_1_sgdma_csr_write,        --                 .write
			csr_writedata                 => mm_interconnect_1_sgdma_csr_writedata,    --                 .writedata
			csr_readdata                  => mm_interconnect_1_sgdma_csr_readdata,     --                 .readdata
			descriptor_read_readdata      => sgdma_descriptor_read_readdata,           --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_descriptor_read_readdatavalid,      --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_descriptor_read_waitrequest,        --                 .waitrequest
			descriptor_read_address       => sgdma_descriptor_read_address,            --                 .address
			descriptor_read_read          => sgdma_descriptor_read_read,               --                 .read
			descriptor_write_waitrequest  => sgdma_descriptor_write_waitrequest,       -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_descriptor_write_address,           --                 .address
			descriptor_write_write        => sgdma_descriptor_write_write,             --                 .write
			descriptor_write_writedata    => sgdma_descriptor_write_writedata,         --                 .writedata
			csr_irq                       => irq_mapper_receiver0_irq,                 --          csr_irq.irq
			m_read_readdata               => sgdma_m_read_readdata,                    --           m_read.readdata
			m_read_readdatavalid          => sgdma_m_read_readdatavalid,               --                 .readdatavalid
			m_read_waitrequest            => sgdma_m_read_waitrequest,                 --                 .waitrequest
			m_read_address                => sgdma_m_read_address,                     --                 .address
			m_read_read                   => sgdma_m_read_read,                        --                 .read
			m_write_waitrequest           => sgdma_m_write_waitrequest,                --          m_write.waitrequest
			m_write_address               => sgdma_m_write_address,                    --                 .address
			m_write_write                 => sgdma_m_write_write,                      --                 .write
			m_write_writedata             => sgdma_m_write_writedata,                  --                 .writedata
			m_write_byteenable            => sgdma_m_write_byteenable                  --                 .byteenable
		);

	fir_memory : component de2i_150_qsys_fir_memory
		port map (
			clk         => pcie_ip_pcie_core_clk_clk,                  --   clk1.clk
			address     => mm_interconnect_0_fir_memory_s1_address,    --     s1.address
			clken       => mm_interconnect_0_fir_memory_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_fir_memory_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_fir_memory_s1_write,      --       .write
			readdata    => mm_interconnect_0_fir_memory_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_fir_memory_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_fir_memory_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,         --       .reset_req
			address2    => fir_memory_s2_address,                      --     s2.address
			chipselect2 => fir_memory_s2_chipselect,                   --       .chipselect
			clken2      => fir_memory_s2_clken,                        --       .clken
			write2      => fir_memory_s2_write,                        --       .write
			readdata2   => fir_memory_s2_readdata,                     --       .readdata
			writedata2  => fir_memory_s2_writedata,                    --       .writedata
			byteenable2 => fir_memory_s2_byteenable,                   --       .byteenable
			clk2        => fir_memory_clk2_clk,                        --   clk2.clk
			reset2      => fir_memory_reset2_reset,                    -- reset2.reset
			reset_req2  => fir_memory_reset2_reset_req                 --       .reset_req
		);

	led : component de2i_150_qsys_led
		port map (
			clk        => pcie_ip_pcie_core_clk_clk,                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,        --                    .readdata
			out_port   => led_external_connection_export            -- external_connection.export
		);

	button : component de2i_150_qsys_button
		port map (
			clk        => pcie_ip_pcie_core_clk_clk,                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_button_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_button_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_button_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_button_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_button_s1_readdata,        --                    .readdata
			in_port    => button_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver2_irq                     --                 irq.irq
		);

	fifo_memory : component de2i_150_qsys_fifo_memory
		port map (
			wrclock                          => pcie_ip_pcie_core_clk_clk,                      --   clk_in.clk
			reset_n                          => rst_controller_reset_out_reset_ports_inv,       -- reset_in.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_0_fifo_memory_in_writedata,     --       in.writedata
			avalonmm_write_slave_write       => mm_interconnect_0_fifo_memory_in_write,         --         .write
			avalonmm_write_slave_waitrequest => mm_interconnect_0_fifo_memory_in_waitrequest,   --         .waitrequest
			avalonmm_read_slave_readdata     => mm_interconnect_0_fifo_memory_out_readdata,     --      out.readdata
			avalonmm_read_slave_read         => mm_interconnect_0_fifo_memory_out_read,         --         .read
			avalonmm_read_slave_waitrequest  => mm_interconnect_0_fifo_memory_out_waitrequest,  --         .waitrequest
			wrclk_control_slave_address      => mm_interconnect_0_fifo_memory_in_csr_address,   --   in_csr.address
			wrclk_control_slave_read         => mm_interconnect_0_fifo_memory_in_csr_read,      --         .read
			wrclk_control_slave_writedata    => mm_interconnect_0_fifo_memory_in_csr_writedata, --         .writedata
			wrclk_control_slave_write        => mm_interconnect_0_fifo_memory_in_csr_write,     --         .write
			wrclk_control_slave_readdata     => mm_interconnect_0_fifo_memory_in_csr_readdata,  --         .readdata
			wrclk_control_slave_irq          => irq_mapper_receiver1_irq                        --   in_irq.irq
		);

	interpo_4_0 : component de2i_150_qsys_Interpo_4_0
		port map (
			clk         => pcie_ip_pcie_core_clk_clk,                   --   clk1.clk
			address     => mm_interconnect_0_interpo_4_0_s1_address,    --     s1.address
			clken       => mm_interconnect_0_interpo_4_0_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_interpo_4_0_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_interpo_4_0_s1_write,      --       .write
			readdata    => mm_interconnect_0_interpo_4_0_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_interpo_4_0_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_interpo_4_0_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,          --       .reset_req
			address2    => interpo_4_0_s2_address,                      --     s2.address
			chipselect2 => interpo_4_0_s2_chipselect,                   --       .chipselect
			clken2      => interpo_4_0_s2_clken,                        --       .clken
			write2      => interpo_4_0_s2_write,                        --       .write
			readdata2   => interpo_4_0_s2_readdata,                     --       .readdata
			writedata2  => interpo_4_0_s2_writedata,                    --       .writedata
			byteenable2 => interpo_4_0_s2_byteenable,                   --       .byteenable
			clk2        => interpo_4_0_clk2_clk,                        --   clk2.clk
			reset2      => interpo_4_0_reset2_reset,                    -- reset2.reset
			reset_req2  => interpo_4_0_reset2_reset_req                 --       .reset_req
		);

	interpo_5_0 : component de2i_150_qsys_Interpo_5_0
		port map (
			clk         => pcie_ip_pcie_core_clk_clk,                   --   clk1.clk
			address     => mm_interconnect_0_interpo_5_0_s1_address,    --     s1.address
			clken       => mm_interconnect_0_interpo_5_0_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_interpo_5_0_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_interpo_5_0_s1_write,      --       .write
			readdata    => mm_interconnect_0_interpo_5_0_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_interpo_5_0_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_interpo_5_0_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,          --       .reset_req
			address2    => interpo_5_0_s2_address,                      --     s2.address
			chipselect2 => interpo_5_0_s2_chipselect,                   --       .chipselect
			clken2      => interpo_5_0_s2_clken,                        --       .clken
			write2      => interpo_5_0_s2_write,                        --       .write
			readdata2   => interpo_5_0_s2_readdata,                     --       .readdata
			writedata2  => interpo_5_0_s2_writedata,                    --       .writedata
			byteenable2 => interpo_5_0_s2_byteenable,                   --       .byteenable
			clk2        => interpo_5_0_clk2_clk,                        --   clk2.clk
			reset2      => interpo_5_0_reset2_reset,                    -- reset2.reset
			reset_req2  => interpo_5_0_reset2_reset_req                 --       .reset_req
		);

	interpo_5_1 : component de2i_150_qsys_Interpo_5_1
		port map (
			clk         => pcie_ip_pcie_core_clk_clk,                   --   clk1.clk
			address     => mm_interconnect_0_interpo_5_1_s1_address,    --     s1.address
			clken       => mm_interconnect_0_interpo_5_1_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_interpo_5_1_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_interpo_5_1_s1_write,      --       .write
			readdata    => mm_interconnect_0_interpo_5_1_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_interpo_5_1_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_interpo_5_1_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,          --       .reset_req
			address2    => interpo_5_1_s2_address,                      --     s2.address
			chipselect2 => interpo_5_1_s2_chipselect,                   --       .chipselect
			clken2      => interpo_5_1_s2_clken,                        --       .clken
			write2      => interpo_5_1_s2_write,                        --       .write
			readdata2   => interpo_5_1_s2_readdata,                     --       .readdata
			writedata2  => interpo_5_1_s2_writedata,                    --       .writedata
			byteenable2 => interpo_5_1_s2_byteenable,                   --       .byteenable
			clk2        => interpo_5_1_clk2_clk,                        --   clk2.clk
			reset2      => interpo_5_1_reset2_reset,                    -- reset2.reset
			reset_req2  => interpo_5_1_reset2_reset_req                 --       .reset_req
		);

	interpo_5_2 : component de2i_150_qsys_Interpo_5_2
		port map (
			clk         => pcie_ip_pcie_core_clk_clk,                   --   clk1.clk
			address     => mm_interconnect_0_interpo_5_2_s1_address,    --     s1.address
			clken       => mm_interconnect_0_interpo_5_2_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_interpo_5_2_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_interpo_5_2_s1_write,      --       .write
			readdata    => mm_interconnect_0_interpo_5_2_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_interpo_5_2_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_interpo_5_2_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,          --       .reset_req
			address2    => interpo_5_2_s2_address,                      --     s2.address
			chipselect2 => interpo_5_2_s2_chipselect,                   --       .chipselect
			clken2      => interpo_5_2_s2_clken,                        --       .clken
			write2      => interpo_5_2_s2_write,                        --       .write
			readdata2   => interpo_5_2_s2_readdata,                     --       .readdata
			writedata2  => interpo_5_2_s2_writedata,                    --       .writedata
			byteenable2 => interpo_5_2_s2_byteenable,                   --       .byteenable
			clk2        => interpo_5_2_clk2_clk,                        --   clk2.clk
			reset2      => interpo_5_2_reset2_reset,                    -- reset2.reset
			reset_req2  => interpo_5_2_reset2_reset_req                 --       .reset_req
		);

	interpo_5_3 : component de2i_150_qsys_Interpo_5_3
		port map (
			clk         => pcie_ip_pcie_core_clk_clk,                   --   clk1.clk
			address     => mm_interconnect_0_interpo_5_3_s1_address,    --     s1.address
			clken       => mm_interconnect_0_interpo_5_3_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_interpo_5_3_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_interpo_5_3_s1_write,      --       .write
			readdata    => mm_interconnect_0_interpo_5_3_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_interpo_5_3_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_interpo_5_3_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,          --       .reset_req
			address2    => interpo_5_3_s2_address,                      --     s2.address
			chipselect2 => interpo_5_3_s2_chipselect,                   --       .chipselect
			clken2      => interpo_5_3_s2_clken,                        --       .clken
			write2      => interpo_5_3_s2_write,                        --       .write
			readdata2   => interpo_5_3_s2_readdata,                     --       .readdata
			writedata2  => interpo_5_3_s2_writedata,                    --       .writedata
			byteenable2 => interpo_5_3_s2_byteenable,                   --       .byteenable
			clk2        => interpo_5_3_clk2_clk,                        --   clk2.clk
			reset2      => interpo_5_3_reset2_reset,                    -- reset2.reset
			reset_req2  => interpo_5_3_reset2_reset_req                 --       .reset_req
		);

	adapt_fir_mem : component de2i_150_qsys_Adapt_FIR_mem
		port map (
			clk         => pcie_ip_pcie_core_clk_clk,                     --   clk1.clk
			address     => mm_interconnect_0_adapt_fir_mem_s1_address,    --     s1.address
			clken       => mm_interconnect_0_adapt_fir_mem_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_adapt_fir_mem_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_adapt_fir_mem_s1_write,      --       .write
			readdata    => mm_interconnect_0_adapt_fir_mem_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_adapt_fir_mem_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_adapt_fir_mem_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,                -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,            --       .reset_req
			address2    => adapt_fir_mem_s2_address,                      --     s2.address
			chipselect2 => adapt_fir_mem_s2_chipselect,                   --       .chipselect
			clken2      => adapt_fir_mem_s2_clken,                        --       .clken
			write2      => adapt_fir_mem_s2_write,                        --       .write
			readdata2   => adapt_fir_mem_s2_readdata,                     --       .readdata
			writedata2  => adapt_fir_mem_s2_writedata,                    --       .writedata
			byteenable2 => adapt_fir_mem_s2_byteenable,                   --       .byteenable
			clk2        => adapt_fir_mem_clk2_clk,                        --   clk2.clk
			reset2      => adapt_fir_mem_reset2_reset,                    -- reset2.reset
			reset_req2  => adapt_fir_mem_reset2_reset_req                 --       .reset_req
		);

	micfilter_cntl : component de2i_150_qsys_micFilter_cntl
		port map (
			clk        => pcie_ip_pcie_core_clk_clk,                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address    => mm_interconnect_0_micfilter_cntl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_micfilter_cntl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_micfilter_cntl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_micfilter_cntl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_micfilter_cntl_s1_readdata,        --                    .readdata
			out_port   => micfilter_cntl_export                                -- external_connection.export
		);

	micfilter_rst : component de2i_150_qsys_micFilter_rst
		port map (
			clk        => pcie_ip_pcie_core_clk_clk,                          --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address    => mm_interconnect_0_micfilter_rst_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_micfilter_rst_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_micfilter_rst_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_micfilter_rst_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_micfilter_rst_s1_readdata,        --                    .readdata
			out_port   => micfilter_rst_export                                -- external_connection.export
		);

	micfilter_adjust : component de2i_150_qsys_micFilter_rst
		port map (
			clk        => pcie_ip_pcie_core_clk_clk,                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_0_micfilter_adjust_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_micfilter_adjust_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_micfilter_adjust_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_micfilter_adjust_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_micfilter_adjust_s1_readdata,        --                    .readdata
			out_port   => micfilter_adjust_export                                -- external_connection.export
		);

	mm_interconnect_0 : component de2i_150_qsys_mm_interconnect_0
		port map (
			pcie_ip_pcie_core_clk_clk                                   => pcie_ip_pcie_core_clk_clk,                        --                                 pcie_ip_pcie_core_clk.clk
			pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,               -- pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset.reset
			sgdma_reset_reset_bridge_in_reset_reset                     => rst_controller_reset_out_reset,                   --                     sgdma_reset_reset_bridge_in_reset.reset
			pcie_ip_bar1_0_address                                      => pcie_ip_bar1_0_address,                           --                                        pcie_ip_bar1_0.address
			pcie_ip_bar1_0_waitrequest                                  => pcie_ip_bar1_0_waitrequest,                       --                                                      .waitrequest
			pcie_ip_bar1_0_burstcount                                   => pcie_ip_bar1_0_burstcount,                        --                                                      .burstcount
			pcie_ip_bar1_0_byteenable                                   => pcie_ip_bar1_0_byteenable,                        --                                                      .byteenable
			pcie_ip_bar1_0_read                                         => pcie_ip_bar1_0_read,                              --                                                      .read
			pcie_ip_bar1_0_readdata                                     => pcie_ip_bar1_0_readdata,                          --                                                      .readdata
			pcie_ip_bar1_0_readdatavalid                                => pcie_ip_bar1_0_readdatavalid,                     --                                                      .readdatavalid
			pcie_ip_bar1_0_write                                        => pcie_ip_bar1_0_write,                             --                                                      .write
			pcie_ip_bar1_0_writedata                                    => pcie_ip_bar1_0_writedata,                         --                                                      .writedata
			sgdma_descriptor_read_address                               => sgdma_descriptor_read_address,                    --                                 sgdma_descriptor_read.address
			sgdma_descriptor_read_waitrequest                           => sgdma_descriptor_read_waitrequest,                --                                                      .waitrequest
			sgdma_descriptor_read_read                                  => sgdma_descriptor_read_read,                       --                                                      .read
			sgdma_descriptor_read_readdata                              => sgdma_descriptor_read_readdata,                   --                                                      .readdata
			sgdma_descriptor_read_readdatavalid                         => sgdma_descriptor_read_readdatavalid,              --                                                      .readdatavalid
			sgdma_descriptor_write_address                              => sgdma_descriptor_write_address,                   --                                sgdma_descriptor_write.address
			sgdma_descriptor_write_waitrequest                          => sgdma_descriptor_write_waitrequest,               --                                                      .waitrequest
			sgdma_descriptor_write_write                                => sgdma_descriptor_write_write,                     --                                                      .write
			sgdma_descriptor_write_writedata                            => sgdma_descriptor_write_writedata,                 --                                                      .writedata
			sgdma_m_read_address                                        => sgdma_m_read_address,                             --                                          sgdma_m_read.address
			sgdma_m_read_waitrequest                                    => sgdma_m_read_waitrequest,                         --                                                      .waitrequest
			sgdma_m_read_read                                           => sgdma_m_read_read,                                --                                                      .read
			sgdma_m_read_readdata                                       => sgdma_m_read_readdata,                            --                                                      .readdata
			sgdma_m_read_readdatavalid                                  => sgdma_m_read_readdatavalid,                       --                                                      .readdatavalid
			sgdma_m_write_address                                       => sgdma_m_write_address,                            --                                         sgdma_m_write.address
			sgdma_m_write_waitrequest                                   => sgdma_m_write_waitrequest,                        --                                                      .waitrequest
			sgdma_m_write_byteenable                                    => sgdma_m_write_byteenable,                         --                                                      .byteenable
			sgdma_m_write_write                                         => sgdma_m_write_write,                              --                                                      .write
			sgdma_m_write_writedata                                     => sgdma_m_write_writedata,                          --                                                      .writedata
			Adapt_FIR_mem_s1_address                                    => mm_interconnect_0_adapt_fir_mem_s1_address,       --                                      Adapt_FIR_mem_s1.address
			Adapt_FIR_mem_s1_write                                      => mm_interconnect_0_adapt_fir_mem_s1_write,         --                                                      .write
			Adapt_FIR_mem_s1_readdata                                   => mm_interconnect_0_adapt_fir_mem_s1_readdata,      --                                                      .readdata
			Adapt_FIR_mem_s1_writedata                                  => mm_interconnect_0_adapt_fir_mem_s1_writedata,     --                                                      .writedata
			Adapt_FIR_mem_s1_byteenable                                 => mm_interconnect_0_adapt_fir_mem_s1_byteenable,    --                                                      .byteenable
			Adapt_FIR_mem_s1_chipselect                                 => mm_interconnect_0_adapt_fir_mem_s1_chipselect,    --                                                      .chipselect
			Adapt_FIR_mem_s1_clken                                      => mm_interconnect_0_adapt_fir_mem_s1_clken,         --                                                      .clken
			button_s1_address                                           => mm_interconnect_0_button_s1_address,              --                                             button_s1.address
			button_s1_write                                             => mm_interconnect_0_button_s1_write,                --                                                      .write
			button_s1_readdata                                          => mm_interconnect_0_button_s1_readdata,             --                                                      .readdata
			button_s1_writedata                                         => mm_interconnect_0_button_s1_writedata,            --                                                      .writedata
			button_s1_chipselect                                        => mm_interconnect_0_button_s1_chipselect,           --                                                      .chipselect
			fifo_memory_in_write                                        => mm_interconnect_0_fifo_memory_in_write,           --                                        fifo_memory_in.write
			fifo_memory_in_writedata                                    => mm_interconnect_0_fifo_memory_in_writedata,       --                                                      .writedata
			fifo_memory_in_waitrequest                                  => mm_interconnect_0_fifo_memory_in_waitrequest,     --                                                      .waitrequest
			fifo_memory_in_csr_address                                  => mm_interconnect_0_fifo_memory_in_csr_address,     --                                    fifo_memory_in_csr.address
			fifo_memory_in_csr_write                                    => mm_interconnect_0_fifo_memory_in_csr_write,       --                                                      .write
			fifo_memory_in_csr_read                                     => mm_interconnect_0_fifo_memory_in_csr_read,        --                                                      .read
			fifo_memory_in_csr_readdata                                 => mm_interconnect_0_fifo_memory_in_csr_readdata,    --                                                      .readdata
			fifo_memory_in_csr_writedata                                => mm_interconnect_0_fifo_memory_in_csr_writedata,   --                                                      .writedata
			fifo_memory_out_read                                        => mm_interconnect_0_fifo_memory_out_read,           --                                       fifo_memory_out.read
			fifo_memory_out_readdata                                    => mm_interconnect_0_fifo_memory_out_readdata,       --                                                      .readdata
			fifo_memory_out_waitrequest                                 => mm_interconnect_0_fifo_memory_out_waitrequest,    --                                                      .waitrequest
			fir_memory_s1_address                                       => mm_interconnect_0_fir_memory_s1_address,          --                                         fir_memory_s1.address
			fir_memory_s1_write                                         => mm_interconnect_0_fir_memory_s1_write,            --                                                      .write
			fir_memory_s1_readdata                                      => mm_interconnect_0_fir_memory_s1_readdata,         --                                                      .readdata
			fir_memory_s1_writedata                                     => mm_interconnect_0_fir_memory_s1_writedata,        --                                                      .writedata
			fir_memory_s1_byteenable                                    => mm_interconnect_0_fir_memory_s1_byteenable,       --                                                      .byteenable
			fir_memory_s1_chipselect                                    => mm_interconnect_0_fir_memory_s1_chipselect,       --                                                      .chipselect
			fir_memory_s1_clken                                         => mm_interconnect_0_fir_memory_s1_clken,            --                                                      .clken
			Interpo_4_0_s1_address                                      => mm_interconnect_0_interpo_4_0_s1_address,         --                                        Interpo_4_0_s1.address
			Interpo_4_0_s1_write                                        => mm_interconnect_0_interpo_4_0_s1_write,           --                                                      .write
			Interpo_4_0_s1_readdata                                     => mm_interconnect_0_interpo_4_0_s1_readdata,        --                                                      .readdata
			Interpo_4_0_s1_writedata                                    => mm_interconnect_0_interpo_4_0_s1_writedata,       --                                                      .writedata
			Interpo_4_0_s1_byteenable                                   => mm_interconnect_0_interpo_4_0_s1_byteenable,      --                                                      .byteenable
			Interpo_4_0_s1_chipselect                                   => mm_interconnect_0_interpo_4_0_s1_chipselect,      --                                                      .chipselect
			Interpo_4_0_s1_clken                                        => mm_interconnect_0_interpo_4_0_s1_clken,           --                                                      .clken
			Interpo_5_0_s1_address                                      => mm_interconnect_0_interpo_5_0_s1_address,         --                                        Interpo_5_0_s1.address
			Interpo_5_0_s1_write                                        => mm_interconnect_0_interpo_5_0_s1_write,           --                                                      .write
			Interpo_5_0_s1_readdata                                     => mm_interconnect_0_interpo_5_0_s1_readdata,        --                                                      .readdata
			Interpo_5_0_s1_writedata                                    => mm_interconnect_0_interpo_5_0_s1_writedata,       --                                                      .writedata
			Interpo_5_0_s1_byteenable                                   => mm_interconnect_0_interpo_5_0_s1_byteenable,      --                                                      .byteenable
			Interpo_5_0_s1_chipselect                                   => mm_interconnect_0_interpo_5_0_s1_chipselect,      --                                                      .chipselect
			Interpo_5_0_s1_clken                                        => mm_interconnect_0_interpo_5_0_s1_clken,           --                                                      .clken
			Interpo_5_1_s1_address                                      => mm_interconnect_0_interpo_5_1_s1_address,         --                                        Interpo_5_1_s1.address
			Interpo_5_1_s1_write                                        => mm_interconnect_0_interpo_5_1_s1_write,           --                                                      .write
			Interpo_5_1_s1_readdata                                     => mm_interconnect_0_interpo_5_1_s1_readdata,        --                                                      .readdata
			Interpo_5_1_s1_writedata                                    => mm_interconnect_0_interpo_5_1_s1_writedata,       --                                                      .writedata
			Interpo_5_1_s1_byteenable                                   => mm_interconnect_0_interpo_5_1_s1_byteenable,      --                                                      .byteenable
			Interpo_5_1_s1_chipselect                                   => mm_interconnect_0_interpo_5_1_s1_chipselect,      --                                                      .chipselect
			Interpo_5_1_s1_clken                                        => mm_interconnect_0_interpo_5_1_s1_clken,           --                                                      .clken
			Interpo_5_2_s1_address                                      => mm_interconnect_0_interpo_5_2_s1_address,         --                                        Interpo_5_2_s1.address
			Interpo_5_2_s1_write                                        => mm_interconnect_0_interpo_5_2_s1_write,           --                                                      .write
			Interpo_5_2_s1_readdata                                     => mm_interconnect_0_interpo_5_2_s1_readdata,        --                                                      .readdata
			Interpo_5_2_s1_writedata                                    => mm_interconnect_0_interpo_5_2_s1_writedata,       --                                                      .writedata
			Interpo_5_2_s1_byteenable                                   => mm_interconnect_0_interpo_5_2_s1_byteenable,      --                                                      .byteenable
			Interpo_5_2_s1_chipselect                                   => mm_interconnect_0_interpo_5_2_s1_chipselect,      --                                                      .chipselect
			Interpo_5_2_s1_clken                                        => mm_interconnect_0_interpo_5_2_s1_clken,           --                                                      .clken
			Interpo_5_3_s1_address                                      => mm_interconnect_0_interpo_5_3_s1_address,         --                                        Interpo_5_3_s1.address
			Interpo_5_3_s1_write                                        => mm_interconnect_0_interpo_5_3_s1_write,           --                                                      .write
			Interpo_5_3_s1_readdata                                     => mm_interconnect_0_interpo_5_3_s1_readdata,        --                                                      .readdata
			Interpo_5_3_s1_writedata                                    => mm_interconnect_0_interpo_5_3_s1_writedata,       --                                                      .writedata
			Interpo_5_3_s1_byteenable                                   => mm_interconnect_0_interpo_5_3_s1_byteenable,      --                                                      .byteenable
			Interpo_5_3_s1_chipselect                                   => mm_interconnect_0_interpo_5_3_s1_chipselect,      --                                                      .chipselect
			Interpo_5_3_s1_clken                                        => mm_interconnect_0_interpo_5_3_s1_clken,           --                                                      .clken
			led_s1_address                                              => mm_interconnect_0_led_s1_address,                 --                                                led_s1.address
			led_s1_write                                                => mm_interconnect_0_led_s1_write,                   --                                                      .write
			led_s1_readdata                                             => mm_interconnect_0_led_s1_readdata,                --                                                      .readdata
			led_s1_writedata                                            => mm_interconnect_0_led_s1_writedata,               --                                                      .writedata
			led_s1_chipselect                                           => mm_interconnect_0_led_s1_chipselect,              --                                                      .chipselect
			micFilter_adjust_s1_address                                 => mm_interconnect_0_micfilter_adjust_s1_address,    --                                   micFilter_adjust_s1.address
			micFilter_adjust_s1_write                                   => mm_interconnect_0_micfilter_adjust_s1_write,      --                                                      .write
			micFilter_adjust_s1_readdata                                => mm_interconnect_0_micfilter_adjust_s1_readdata,   --                                                      .readdata
			micFilter_adjust_s1_writedata                               => mm_interconnect_0_micfilter_adjust_s1_writedata,  --                                                      .writedata
			micFilter_adjust_s1_chipselect                              => mm_interconnect_0_micfilter_adjust_s1_chipselect, --                                                      .chipselect
			micFilter_cntl_s1_address                                   => mm_interconnect_0_micfilter_cntl_s1_address,      --                                     micFilter_cntl_s1.address
			micFilter_cntl_s1_write                                     => mm_interconnect_0_micfilter_cntl_s1_write,        --                                                      .write
			micFilter_cntl_s1_readdata                                  => mm_interconnect_0_micfilter_cntl_s1_readdata,     --                                                      .readdata
			micFilter_cntl_s1_writedata                                 => mm_interconnect_0_micfilter_cntl_s1_writedata,    --                                                      .writedata
			micFilter_cntl_s1_chipselect                                => mm_interconnect_0_micfilter_cntl_s1_chipselect,   --                                                      .chipselect
			micFilter_rst_s1_address                                    => mm_interconnect_0_micfilter_rst_s1_address,       --                                      micFilter_rst_s1.address
			micFilter_rst_s1_write                                      => mm_interconnect_0_micfilter_rst_s1_write,         --                                                      .write
			micFilter_rst_s1_readdata                                   => mm_interconnect_0_micfilter_rst_s1_readdata,      --                                                      .readdata
			micFilter_rst_s1_writedata                                  => mm_interconnect_0_micfilter_rst_s1_writedata,     --                                                      .writedata
			micFilter_rst_s1_chipselect                                 => mm_interconnect_0_micfilter_rst_s1_chipselect,    --                                                      .chipselect
			pcie_ip_txs_address                                         => mm_interconnect_0_pcie_ip_txs_address,            --                                           pcie_ip_txs.address
			pcie_ip_txs_write                                           => mm_interconnect_0_pcie_ip_txs_write,              --                                                      .write
			pcie_ip_txs_read                                            => mm_interconnect_0_pcie_ip_txs_read,               --                                                      .read
			pcie_ip_txs_readdata                                        => mm_interconnect_0_pcie_ip_txs_readdata,           --                                                      .readdata
			pcie_ip_txs_writedata                                       => mm_interconnect_0_pcie_ip_txs_writedata,          --                                                      .writedata
			pcie_ip_txs_burstcount                                      => mm_interconnect_0_pcie_ip_txs_burstcount,         --                                                      .burstcount
			pcie_ip_txs_byteenable                                      => mm_interconnect_0_pcie_ip_txs_byteenable,         --                                                      .byteenable
			pcie_ip_txs_readdatavalid                                   => mm_interconnect_0_pcie_ip_txs_readdatavalid,      --                                                      .readdatavalid
			pcie_ip_txs_waitrequest                                     => mm_interconnect_0_pcie_ip_txs_waitrequest,        --                                                      .waitrequest
			pcie_ip_txs_chipselect                                      => mm_interconnect_0_pcie_ip_txs_chipselect          --                                                      .chipselect
		);

	mm_interconnect_1 : component de2i_150_qsys_mm_interconnect_1
		port map (
			pcie_ip_pcie_core_clk_clk                                 => pcie_ip_pcie_core_clk_clk,                 --                               pcie_ip_pcie_core_clk.clk
			pcie_ip_bar2_translator_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,        -- pcie_ip_bar2_translator_reset_reset_bridge_in_reset.reset
			sgdma_reset_reset_bridge_in_reset_reset                   => rst_controller_reset_out_reset,            --                   sgdma_reset_reset_bridge_in_reset.reset
			pcie_ip_bar2_address                                      => pcie_ip_bar2_address,                      --                                        pcie_ip_bar2.address
			pcie_ip_bar2_waitrequest                                  => pcie_ip_bar2_waitrequest,                  --                                                    .waitrequest
			pcie_ip_bar2_burstcount                                   => pcie_ip_bar2_burstcount,                   --                                                    .burstcount
			pcie_ip_bar2_byteenable                                   => pcie_ip_bar2_byteenable,                   --                                                    .byteenable
			pcie_ip_bar2_read                                         => pcie_ip_bar2_read,                         --                                                    .read
			pcie_ip_bar2_readdata                                     => pcie_ip_bar2_readdata,                     --                                                    .readdata
			pcie_ip_bar2_readdatavalid                                => pcie_ip_bar2_readdatavalid,                --                                                    .readdatavalid
			pcie_ip_bar2_write                                        => pcie_ip_bar2_write,                        --                                                    .write
			pcie_ip_bar2_writedata                                    => pcie_ip_bar2_writedata,                    --                                                    .writedata
			pcie_ip_cra_address                                       => mm_interconnect_1_pcie_ip_cra_address,     --                                         pcie_ip_cra.address
			pcie_ip_cra_write                                         => mm_interconnect_1_pcie_ip_cra_write,       --                                                    .write
			pcie_ip_cra_read                                          => mm_interconnect_1_pcie_ip_cra_read,        --                                                    .read
			pcie_ip_cra_readdata                                      => mm_interconnect_1_pcie_ip_cra_readdata,    --                                                    .readdata
			pcie_ip_cra_writedata                                     => mm_interconnect_1_pcie_ip_cra_writedata,   --                                                    .writedata
			pcie_ip_cra_byteenable                                    => mm_interconnect_1_pcie_ip_cra_byteenable,  --                                                    .byteenable
			pcie_ip_cra_waitrequest                                   => mm_interconnect_1_pcie_ip_cra_waitrequest, --                                                    .waitrequest
			pcie_ip_cra_chipselect                                    => mm_interconnect_1_pcie_ip_cra_chipselect,  --                                                    .chipselect
			sgdma_csr_address                                         => mm_interconnect_1_sgdma_csr_address,       --                                           sgdma_csr.address
			sgdma_csr_write                                           => mm_interconnect_1_sgdma_csr_write,         --                                                    .write
			sgdma_csr_read                                            => mm_interconnect_1_sgdma_csr_read,          --                                                    .read
			sgdma_csr_readdata                                        => mm_interconnect_1_sgdma_csr_readdata,      --                                                    .readdata
			sgdma_csr_writedata                                       => mm_interconnect_1_sgdma_csr_writedata,     --                                                    .writedata
			sgdma_csr_chipselect                                      => mm_interconnect_1_sgdma_csr_chipselect     --                                                    .chipselect
		);

	irq_mapper : component de2i_150_qsys_irq_mapper
		port map (
			clk           => pcie_ip_pcie_core_clk_clk,          --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			sender_irq    => pcie_ip_rxm_irq_irq                 --    sender.irq
		);

	rst_controller : component de2i_150_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => pcie_ip_pcie_core_reset_reset_ports_inv, -- reset_in0.reset
			reset_in1      => reset_reset_n_ports_inv,                 -- reset_in1.reset
			clk            => pcie_ip_pcie_core_clk_clk,               --       clk.clk
			reset_out      => rst_controller_reset_out_reset,          -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,      --          .reset_req
			reset_req_in0  => '0',                                     -- (terminated)
			reset_req_in1  => '0',                                     -- (terminated)
			reset_in2      => '0',                                     -- (terminated)
			reset_req_in2  => '0',                                     -- (terminated)
			reset_in3      => '0',                                     -- (terminated)
			reset_req_in3  => '0',                                     -- (terminated)
			reset_in4      => '0',                                     -- (terminated)
			reset_req_in4  => '0',                                     -- (terminated)
			reset_in5      => '0',                                     -- (terminated)
			reset_req_in5  => '0',                                     -- (terminated)
			reset_in6      => '0',                                     -- (terminated)
			reset_req_in6  => '0',                                     -- (terminated)
			reset_in7      => '0',                                     -- (terminated)
			reset_req_in7  => '0',                                     -- (terminated)
			reset_in8      => '0',                                     -- (terminated)
			reset_req_in8  => '0',                                     -- (terminated)
			reset_in9      => '0',                                     -- (terminated)
			reset_req_in9  => '0',                                     -- (terminated)
			reset_in10     => '0',                                     -- (terminated)
			reset_req_in10 => '0',                                     -- (terminated)
			reset_in11     => '0',                                     -- (terminated)
			reset_req_in11 => '0',                                     -- (terminated)
			reset_in12     => '0',                                     -- (terminated)
			reset_req_in12 => '0',                                     -- (terminated)
			reset_in13     => '0',                                     -- (terminated)
			reset_req_in13 => '0',                                     -- (terminated)
			reset_in14     => '0',                                     -- (terminated)
			reset_req_in14 => '0',                                     -- (terminated)
			reset_in15     => '0',                                     -- (terminated)
			reset_req_in15 => '0'                                      -- (terminated)
		);

	rst_controller_001 : component de2i_150_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => pcie_ip_pcie_core_reset_reset_ports_inv, -- reset_in0.reset
			clk            => pcie_ip_pcie_core_clk_clk,               --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,      -- reset_out.reset
			reset_req      => open,                                    -- (terminated)
			reset_req_in0  => '0',                                     -- (terminated)
			reset_in1      => '0',                                     -- (terminated)
			reset_req_in1  => '0',                                     -- (terminated)
			reset_in2      => '0',                                     -- (terminated)
			reset_req_in2  => '0',                                     -- (terminated)
			reset_in3      => '0',                                     -- (terminated)
			reset_req_in3  => '0',                                     -- (terminated)
			reset_in4      => '0',                                     -- (terminated)
			reset_req_in4  => '0',                                     -- (terminated)
			reset_in5      => '0',                                     -- (terminated)
			reset_req_in5  => '0',                                     -- (terminated)
			reset_in6      => '0',                                     -- (terminated)
			reset_req_in6  => '0',                                     -- (terminated)
			reset_in7      => '0',                                     -- (terminated)
			reset_req_in7  => '0',                                     -- (terminated)
			reset_in8      => '0',                                     -- (terminated)
			reset_req_in8  => '0',                                     -- (terminated)
			reset_in9      => '0',                                     -- (terminated)
			reset_req_in9  => '0',                                     -- (terminated)
			reset_in10     => '0',                                     -- (terminated)
			reset_req_in10 => '0',                                     -- (terminated)
			reset_in11     => '0',                                     -- (terminated)
			reset_req_in11 => '0',                                     -- (terminated)
			reset_in12     => '0',                                     -- (terminated)
			reset_req_in12 => '0',                                     -- (terminated)
			reset_in13     => '0',                                     -- (terminated)
			reset_req_in13 => '0',                                     -- (terminated)
			reset_in14     => '0',                                     -- (terminated)
			reset_req_in14 => '0',                                     -- (terminated)
			reset_in15     => '0',                                     -- (terminated)
			reset_req_in15 => '0'                                      -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	mm_interconnect_0_button_s1_write_ports_inv <= not mm_interconnect_0_button_s1_write;

	mm_interconnect_0_micfilter_cntl_s1_write_ports_inv <= not mm_interconnect_0_micfilter_cntl_s1_write;

	mm_interconnect_0_micfilter_rst_s1_write_ports_inv <= not mm_interconnect_0_micfilter_rst_s1_write;

	mm_interconnect_0_micfilter_adjust_s1_write_ports_inv <= not mm_interconnect_0_micfilter_adjust_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	pcie_ip_pcie_core_reset_reset_ports_inv <= not pcie_ip_pcie_core_reset_reset;

end architecture rtl; -- of de2i_150_qsys
