// de2i_150_qsys.v

// Generated using ACDS version 14.0 200 at 2015.11.29.16:33:49

`timescale 1 ps / 1 ps
module de2i_150_qsys (
		input  wire        clk_clk,                                    //                        clk.clk
		input  wire        reset_reset_n,                              //                      reset.reset_n
		input  wire [3:0]  pcie_ip_reconfig_togxb_data,                //     pcie_ip_reconfig_togxb.data
		input  wire        pcie_ip_refclk_export,                      //             pcie_ip_refclk.export
		input  wire [39:0] pcie_ip_test_in_test_in,                    //            pcie_ip_test_in.test_in
		input  wire        pcie_ip_pcie_rstn_export,                   //          pcie_ip_pcie_rstn.export
		output wire        pcie_ip_clocks_sim_clk250_export,           //         pcie_ip_clocks_sim.clk250_export
		output wire        pcie_ip_clocks_sim_clk500_export,           //                           .clk500_export
		output wire        pcie_ip_clocks_sim_clk125_export,           //                           .clk125_export
		input  wire        pcie_ip_reconfig_busy_busy_altgxb_reconfig, //      pcie_ip_reconfig_busy.busy_altgxb_reconfig
		input  wire        pcie_ip_pipe_ext_pipe_mode,                 //           pcie_ip_pipe_ext.pipe_mode
		input  wire        pcie_ip_pipe_ext_phystatus_ext,             //                           .phystatus_ext
		output wire        pcie_ip_pipe_ext_rate_ext,                  //                           .rate_ext
		output wire [1:0]  pcie_ip_pipe_ext_powerdown_ext,             //                           .powerdown_ext
		output wire        pcie_ip_pipe_ext_txdetectrx_ext,            //                           .txdetectrx_ext
		input  wire        pcie_ip_pipe_ext_rxelecidle0_ext,           //                           .rxelecidle0_ext
		input  wire [7:0]  pcie_ip_pipe_ext_rxdata0_ext,               //                           .rxdata0_ext
		input  wire [2:0]  pcie_ip_pipe_ext_rxstatus0_ext,             //                           .rxstatus0_ext
		input  wire        pcie_ip_pipe_ext_rxvalid0_ext,              //                           .rxvalid0_ext
		input  wire        pcie_ip_pipe_ext_rxdatak0_ext,              //                           .rxdatak0_ext
		output wire [7:0]  pcie_ip_pipe_ext_txdata0_ext,               //                           .txdata0_ext
		output wire        pcie_ip_pipe_ext_txdatak0_ext,              //                           .txdatak0_ext
		output wire        pcie_ip_pipe_ext_rxpolarity0_ext,           //                           .rxpolarity0_ext
		output wire        pcie_ip_pipe_ext_txcompl0_ext,              //                           .txcompl0_ext
		output wire        pcie_ip_pipe_ext_txelecidle0_ext,           //                           .txelecidle0_ext
		input  wire        pcie_ip_rx_in_rx_datain_0,                  //              pcie_ip_rx_in.rx_datain_0
		output wire        pcie_ip_tx_out_tx_dataout_0,                //             pcie_ip_tx_out.tx_dataout_0
		output wire [4:0]  pcie_ip_reconfig_fromgxb_0_data,            // pcie_ip_reconfig_fromgxb_0.data
		output wire [3:0]  led_external_connection_export,             //    led_external_connection.export
		input  wire [3:0]  button_external_connection_export,          // button_external_connection.export
		input  wire [9:0]  fir_memory_s2_address,                      //              fir_memory_s2.address
		input  wire        fir_memory_s2_chipselect,                   //                           .chipselect
		input  wire        fir_memory_s2_clken,                        //                           .clken
		input  wire        fir_memory_s2_write,                        //                           .write
		output wire [31:0] fir_memory_s2_readdata,                     //                           .readdata
		input  wire [31:0] fir_memory_s2_writedata,                    //                           .writedata
		input  wire [3:0]  fir_memory_s2_byteenable,                   //                           .byteenable
		input  wire        fir_memory_clk2_clk,                        //            fir_memory_clk2.clk
		input  wire        fir_memory_reset2_reset,                    //          fir_memory_reset2.reset
		input  wire        fir_memory_reset2_reset_req,                //                           .reset_req
		input  wire [4:0]  interpo_4_0_s2_address,                     //             interpo_4_0_s2.address
		input  wire        interpo_4_0_s2_chipselect,                  //                           .chipselect
		input  wire        interpo_4_0_s2_clken,                       //                           .clken
		input  wire        interpo_4_0_s2_write,                       //                           .write
		output wire [31:0] interpo_4_0_s2_readdata,                    //                           .readdata
		input  wire [31:0] interpo_4_0_s2_writedata,                   //                           .writedata
		input  wire [3:0]  interpo_4_0_s2_byteenable,                  //                           .byteenable
		input  wire        interpo_4_0_clk2_clk,                       //           interpo_4_0_clk2.clk
		input  wire        interpo_4_0_reset2_reset,                   //         interpo_4_0_reset2.reset
		input  wire        interpo_4_0_reset2_reset_req,               //                           .reset_req
		input  wire [5:0]  interpo_5_0_s2_address,                     //             interpo_5_0_s2.address
		input  wire        interpo_5_0_s2_chipselect,                  //                           .chipselect
		input  wire        interpo_5_0_s2_clken,                       //                           .clken
		input  wire        interpo_5_0_s2_write,                       //                           .write
		output wire [31:0] interpo_5_0_s2_readdata,                    //                           .readdata
		input  wire [31:0] interpo_5_0_s2_writedata,                   //                           .writedata
		input  wire [3:0]  interpo_5_0_s2_byteenable,                  //                           .byteenable
		input  wire        interpo_5_0_clk2_clk,                       //           interpo_5_0_clk2.clk
		input  wire        interpo_5_0_reset2_reset,                   //         interpo_5_0_reset2.reset
		input  wire        interpo_5_0_reset2_reset_req,               //                           .reset_req
		input  wire        interpo_5_1_clk2_clk,                       //           interpo_5_1_clk2.clk
		input  wire [5:0]  interpo_5_1_s2_address,                     //             interpo_5_1_s2.address
		input  wire        interpo_5_1_s2_chipselect,                  //                           .chipselect
		input  wire        interpo_5_1_s2_clken,                       //                           .clken
		input  wire        interpo_5_1_s2_write,                       //                           .write
		output wire [31:0] interpo_5_1_s2_readdata,                    //                           .readdata
		input  wire [31:0] interpo_5_1_s2_writedata,                   //                           .writedata
		input  wire [3:0]  interpo_5_1_s2_byteenable,                  //                           .byteenable
		input  wire        interpo_5_1_reset2_reset,                   //         interpo_5_1_reset2.reset
		input  wire        interpo_5_1_reset2_reset_req,               //                           .reset_req
		input  wire [5:0]  interpo_5_2_s2_address,                     //             interpo_5_2_s2.address
		input  wire        interpo_5_2_s2_chipselect,                  //                           .chipselect
		input  wire        interpo_5_2_s2_clken,                       //                           .clken
		input  wire        interpo_5_2_s2_write,                       //                           .write
		output wire [31:0] interpo_5_2_s2_readdata,                    //                           .readdata
		input  wire [31:0] interpo_5_2_s2_writedata,                   //                           .writedata
		input  wire [3:0]  interpo_5_2_s2_byteenable,                  //                           .byteenable
		input  wire        interpo_5_2_clk2_clk,                       //           interpo_5_2_clk2.clk
		input  wire        interpo_5_2_reset2_reset,                   //         interpo_5_2_reset2.reset
		input  wire        interpo_5_2_reset2_reset_req,               //                           .reset_req
		input  wire [5:0]  interpo_5_3_s2_address,                     //             interpo_5_3_s2.address
		input  wire        interpo_5_3_s2_chipselect,                  //                           .chipselect
		input  wire        interpo_5_3_s2_clken,                       //                           .clken
		input  wire        interpo_5_3_s2_write,                       //                           .write
		output wire [31:0] interpo_5_3_s2_readdata,                    //                           .readdata
		input  wire [31:0] interpo_5_3_s2_writedata,                   //                           .writedata
		input  wire [3:0]  interpo_5_3_s2_byteenable,                  //                           .byteenable
		input  wire        interpo_5_3_clk2_clk,                       //           interpo_5_3_clk2.clk
		input  wire        interpo_5_3_reset2_reset,                   //         interpo_5_3_reset2.reset
		input  wire        interpo_5_3_reset2_reset_req,               //                           .reset_req
		input  wire [8:0]  adapt_fir_mem_s2_address,                   //           adapt_fir_mem_s2.address
		input  wire        adapt_fir_mem_s2_chipselect,                //                           .chipselect
		input  wire        adapt_fir_mem_s2_clken,                     //                           .clken
		input  wire        adapt_fir_mem_s2_write,                     //                           .write
		output wire [31:0] adapt_fir_mem_s2_readdata,                  //                           .readdata
		input  wire [31:0] adapt_fir_mem_s2_writedata,                 //                           .writedata
		input  wire [3:0]  adapt_fir_mem_s2_byteenable,                //                           .byteenable
		input  wire        adapt_fir_mem_clk2_clk,                     //         adapt_fir_mem_clk2.clk
		input  wire        adapt_fir_mem_reset2_reset,                 //       adapt_fir_mem_reset2.reset
		input  wire        adapt_fir_mem_reset2_reset_req,             //                           .reset_req
		output wire [31:0] micfilter_cntl_export,                      //             micfilter_cntl.export
		output wire        micfilter_rst_export,                       //              micfilter_rst.export
		output wire        micfilter_adjust_export,                    //           micfilter_adjust.export
		output wire [3:0]  output1_sel_export,                         //                output1_sel.export
		output wire [3:0]  output2_sel_export,                         //                output2_sel.export
		output wire [2:0]  bypass_sel_export,                          //                 bypass_sel.export
		output wire [15:0] sub_factor_export,                          //                 sub_factor.export
		output wire [18:0] delay_lenght_export,                        //               delay_lenght.export
		output wire [31:0] downsamplemult_export,                      //             downsamplemult.export
		output wire [31:0] adapt_weight_export,                        //               adapt_weight.export
		output wire [15:0] adapt_pth_export,                           //                  adapt_pth.export
		output wire [15:0] adapt_nth_export                            //                  adapt_nth.export
	);

	wire         pcie_ip_pcie_core_clk_clk;                        // pcie_ip:pcie_core_clk_clk -> [Adapt_FIR_mem:clk, DownSampleMult:clk, Interpo_4_0:clk, Interpo_5_0:clk, Interpo_5_1:clk, Interpo_5_2:clk, Interpo_5_3:clk, adapt_nTh:clk, adapt_pTh:clk, adapt_weight:clk, button:clk, bypass_sel:clk, delay_lenght:clk, fifo_memory:wrclock, fir_memory:clk, irq_mapper:clk, led:clk, micFilter_adjust:clk, micFilter_cntl:clk, micFilter_rst:clk, mm_interconnect_0:pcie_ip_pcie_core_clk_clk, mm_interconnect_1:pcie_ip_pcie_core_clk_clk, output1_sel:clk, output2_sel:clk, pcie_ip:fixedclk_clk, rst_controller:clk, rst_controller_001:clk, sgdma:clk, sub_factor:clk]
	wire   [6:0] pcie_ip_bar1_0_burstcount;                        // pcie_ip:bar1_0_burstcount -> mm_interconnect_0:pcie_ip_bar1_0_burstcount
	wire         pcie_ip_bar1_0_waitrequest;                       // mm_interconnect_0:pcie_ip_bar1_0_waitrequest -> pcie_ip:bar1_0_waitrequest
	wire  [63:0] pcie_ip_bar1_0_writedata;                         // pcie_ip:bar1_0_writedata -> mm_interconnect_0:pcie_ip_bar1_0_writedata
	wire  [31:0] pcie_ip_bar1_0_address;                           // pcie_ip:bar1_0_address -> mm_interconnect_0:pcie_ip_bar1_0_address
	wire         pcie_ip_bar1_0_write;                             // pcie_ip:bar1_0_write -> mm_interconnect_0:pcie_ip_bar1_0_write
	wire         pcie_ip_bar1_0_read;                              // pcie_ip:bar1_0_read -> mm_interconnect_0:pcie_ip_bar1_0_read
	wire  [63:0] pcie_ip_bar1_0_readdata;                          // mm_interconnect_0:pcie_ip_bar1_0_readdata -> pcie_ip:bar1_0_readdata
	wire   [7:0] pcie_ip_bar1_0_byteenable;                        // pcie_ip:bar1_0_byteenable -> mm_interconnect_0:pcie_ip_bar1_0_byteenable
	wire         pcie_ip_bar1_0_readdatavalid;                     // mm_interconnect_0:pcie_ip_bar1_0_readdatavalid -> pcie_ip:bar1_0_readdatavalid
	wire         sgdma_m_read_waitrequest;                         // mm_interconnect_0:sgdma_m_read_waitrequest -> sgdma:m_read_waitrequest
	wire  [31:0] sgdma_m_read_address;                             // sgdma:m_read_address -> mm_interconnect_0:sgdma_m_read_address
	wire         sgdma_m_read_read;                                // sgdma:m_read_read -> mm_interconnect_0:sgdma_m_read_read
	wire  [63:0] sgdma_m_read_readdata;                            // mm_interconnect_0:sgdma_m_read_readdata -> sgdma:m_read_readdata
	wire         sgdma_m_read_readdatavalid;                       // mm_interconnect_0:sgdma_m_read_readdatavalid -> sgdma:m_read_readdatavalid
	wire         sgdma_m_write_waitrequest;                        // mm_interconnect_0:sgdma_m_write_waitrequest -> sgdma:m_write_waitrequest
	wire  [63:0] sgdma_m_write_writedata;                          // sgdma:m_write_writedata -> mm_interconnect_0:sgdma_m_write_writedata
	wire  [31:0] sgdma_m_write_address;                            // sgdma:m_write_address -> mm_interconnect_0:sgdma_m_write_address
	wire         sgdma_m_write_write;                              // sgdma:m_write_write -> mm_interconnect_0:sgdma_m_write_write
	wire   [7:0] sgdma_m_write_byteenable;                         // sgdma:m_write_byteenable -> mm_interconnect_0:sgdma_m_write_byteenable
	wire         sgdma_descriptor_read_waitrequest;                // mm_interconnect_0:sgdma_descriptor_read_waitrequest -> sgdma:descriptor_read_waitrequest
	wire  [31:0] sgdma_descriptor_read_address;                    // sgdma:descriptor_read_address -> mm_interconnect_0:sgdma_descriptor_read_address
	wire         sgdma_descriptor_read_read;                       // sgdma:descriptor_read_read -> mm_interconnect_0:sgdma_descriptor_read_read
	wire  [31:0] sgdma_descriptor_read_readdata;                   // mm_interconnect_0:sgdma_descriptor_read_readdata -> sgdma:descriptor_read_readdata
	wire         sgdma_descriptor_read_readdatavalid;              // mm_interconnect_0:sgdma_descriptor_read_readdatavalid -> sgdma:descriptor_read_readdatavalid
	wire         sgdma_descriptor_write_waitrequest;               // mm_interconnect_0:sgdma_descriptor_write_waitrequest -> sgdma:descriptor_write_waitrequest
	wire  [31:0] sgdma_descriptor_write_writedata;                 // sgdma:descriptor_write_writedata -> mm_interconnect_0:sgdma_descriptor_write_writedata
	wire  [31:0] sgdma_descriptor_write_address;                   // sgdma:descriptor_write_address -> mm_interconnect_0:sgdma_descriptor_write_address
	wire         sgdma_descriptor_write_write;                     // sgdma:descriptor_write_write -> mm_interconnect_0:sgdma_descriptor_write_write
	wire  [31:0] mm_interconnect_0_fir_memory_s1_writedata;        // mm_interconnect_0:fir_memory_s1_writedata -> fir_memory:writedata
	wire   [9:0] mm_interconnect_0_fir_memory_s1_address;          // mm_interconnect_0:fir_memory_s1_address -> fir_memory:address
	wire         mm_interconnect_0_fir_memory_s1_chipselect;       // mm_interconnect_0:fir_memory_s1_chipselect -> fir_memory:chipselect
	wire         mm_interconnect_0_fir_memory_s1_clken;            // mm_interconnect_0:fir_memory_s1_clken -> fir_memory:clken
	wire         mm_interconnect_0_fir_memory_s1_write;            // mm_interconnect_0:fir_memory_s1_write -> fir_memory:write
	wire  [31:0] mm_interconnect_0_fir_memory_s1_readdata;         // fir_memory:readdata -> mm_interconnect_0:fir_memory_s1_readdata
	wire   [3:0] mm_interconnect_0_fir_memory_s1_byteenable;       // mm_interconnect_0:fir_memory_s1_byteenable -> fir_memory:byteenable
	wire  [31:0] mm_interconnect_0_led_s1_writedata;               // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire   [1:0] mm_interconnect_0_led_s1_address;                 // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_chipselect;              // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire         mm_interconnect_0_led_s1_write;                   // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire  [31:0] mm_interconnect_0_button_s1_writedata;            // mm_interconnect_0:button_s1_writedata -> button:writedata
	wire   [1:0] mm_interconnect_0_button_s1_address;              // mm_interconnect_0:button_s1_address -> button:address
	wire         mm_interconnect_0_button_s1_chipselect;           // mm_interconnect_0:button_s1_chipselect -> button:chipselect
	wire         mm_interconnect_0_button_s1_write;                // mm_interconnect_0:button_s1_write -> button:write_n
	wire  [31:0] mm_interconnect_0_button_s1_readdata;             // button:readdata -> mm_interconnect_0:button_s1_readdata
	wire  [31:0] mm_interconnect_0_fifo_memory_in_csr_writedata;   // mm_interconnect_0:fifo_memory_in_csr_writedata -> fifo_memory:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_memory_in_csr_address;     // mm_interconnect_0:fifo_memory_in_csr_address -> fifo_memory:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_memory_in_csr_write;       // mm_interconnect_0:fifo_memory_in_csr_write -> fifo_memory:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_memory_in_csr_read;        // mm_interconnect_0:fifo_memory_in_csr_read -> fifo_memory:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_memory_in_csr_readdata;    // fifo_memory:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_memory_in_csr_readdata
	wire         mm_interconnect_0_fifo_memory_in_waitrequest;     // fifo_memory:avalonmm_write_slave_waitrequest -> mm_interconnect_0:fifo_memory_in_waitrequest
	wire  [63:0] mm_interconnect_0_fifo_memory_in_writedata;       // mm_interconnect_0:fifo_memory_in_writedata -> fifo_memory:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_memory_in_write;           // mm_interconnect_0:fifo_memory_in_write -> fifo_memory:avalonmm_write_slave_write
	wire         mm_interconnect_0_fifo_memory_out_waitrequest;    // fifo_memory:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_memory_out_waitrequest
	wire         mm_interconnect_0_fifo_memory_out_read;           // mm_interconnect_0:fifo_memory_out_read -> fifo_memory:avalonmm_read_slave_read
	wire  [63:0] mm_interconnect_0_fifo_memory_out_readdata;       // fifo_memory:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_memory_out_readdata
	wire  [31:0] mm_interconnect_0_interpo_4_0_s1_writedata;       // mm_interconnect_0:Interpo_4_0_s1_writedata -> Interpo_4_0:writedata
	wire   [4:0] mm_interconnect_0_interpo_4_0_s1_address;         // mm_interconnect_0:Interpo_4_0_s1_address -> Interpo_4_0:address
	wire         mm_interconnect_0_interpo_4_0_s1_chipselect;      // mm_interconnect_0:Interpo_4_0_s1_chipselect -> Interpo_4_0:chipselect
	wire         mm_interconnect_0_interpo_4_0_s1_clken;           // mm_interconnect_0:Interpo_4_0_s1_clken -> Interpo_4_0:clken
	wire         mm_interconnect_0_interpo_4_0_s1_write;           // mm_interconnect_0:Interpo_4_0_s1_write -> Interpo_4_0:write
	wire  [31:0] mm_interconnect_0_interpo_4_0_s1_readdata;        // Interpo_4_0:readdata -> mm_interconnect_0:Interpo_4_0_s1_readdata
	wire   [3:0] mm_interconnect_0_interpo_4_0_s1_byteenable;      // mm_interconnect_0:Interpo_4_0_s1_byteenable -> Interpo_4_0:byteenable
	wire  [31:0] mm_interconnect_0_interpo_5_0_s1_writedata;       // mm_interconnect_0:Interpo_5_0_s1_writedata -> Interpo_5_0:writedata
	wire   [5:0] mm_interconnect_0_interpo_5_0_s1_address;         // mm_interconnect_0:Interpo_5_0_s1_address -> Interpo_5_0:address
	wire         mm_interconnect_0_interpo_5_0_s1_chipselect;      // mm_interconnect_0:Interpo_5_0_s1_chipselect -> Interpo_5_0:chipselect
	wire         mm_interconnect_0_interpo_5_0_s1_clken;           // mm_interconnect_0:Interpo_5_0_s1_clken -> Interpo_5_0:clken
	wire         mm_interconnect_0_interpo_5_0_s1_write;           // mm_interconnect_0:Interpo_5_0_s1_write -> Interpo_5_0:write
	wire  [31:0] mm_interconnect_0_interpo_5_0_s1_readdata;        // Interpo_5_0:readdata -> mm_interconnect_0:Interpo_5_0_s1_readdata
	wire   [3:0] mm_interconnect_0_interpo_5_0_s1_byteenable;      // mm_interconnect_0:Interpo_5_0_s1_byteenable -> Interpo_5_0:byteenable
	wire  [31:0] mm_interconnect_0_interpo_5_1_s1_writedata;       // mm_interconnect_0:Interpo_5_1_s1_writedata -> Interpo_5_1:writedata
	wire   [5:0] mm_interconnect_0_interpo_5_1_s1_address;         // mm_interconnect_0:Interpo_5_1_s1_address -> Interpo_5_1:address
	wire         mm_interconnect_0_interpo_5_1_s1_chipselect;      // mm_interconnect_0:Interpo_5_1_s1_chipselect -> Interpo_5_1:chipselect
	wire         mm_interconnect_0_interpo_5_1_s1_clken;           // mm_interconnect_0:Interpo_5_1_s1_clken -> Interpo_5_1:clken
	wire         mm_interconnect_0_interpo_5_1_s1_write;           // mm_interconnect_0:Interpo_5_1_s1_write -> Interpo_5_1:write
	wire  [31:0] mm_interconnect_0_interpo_5_1_s1_readdata;        // Interpo_5_1:readdata -> mm_interconnect_0:Interpo_5_1_s1_readdata
	wire   [3:0] mm_interconnect_0_interpo_5_1_s1_byteenable;      // mm_interconnect_0:Interpo_5_1_s1_byteenable -> Interpo_5_1:byteenable
	wire  [31:0] mm_interconnect_0_interpo_5_2_s1_writedata;       // mm_interconnect_0:Interpo_5_2_s1_writedata -> Interpo_5_2:writedata
	wire   [5:0] mm_interconnect_0_interpo_5_2_s1_address;         // mm_interconnect_0:Interpo_5_2_s1_address -> Interpo_5_2:address
	wire         mm_interconnect_0_interpo_5_2_s1_chipselect;      // mm_interconnect_0:Interpo_5_2_s1_chipselect -> Interpo_5_2:chipselect
	wire         mm_interconnect_0_interpo_5_2_s1_clken;           // mm_interconnect_0:Interpo_5_2_s1_clken -> Interpo_5_2:clken
	wire         mm_interconnect_0_interpo_5_2_s1_write;           // mm_interconnect_0:Interpo_5_2_s1_write -> Interpo_5_2:write
	wire  [31:0] mm_interconnect_0_interpo_5_2_s1_readdata;        // Interpo_5_2:readdata -> mm_interconnect_0:Interpo_5_2_s1_readdata
	wire   [3:0] mm_interconnect_0_interpo_5_2_s1_byteenable;      // mm_interconnect_0:Interpo_5_2_s1_byteenable -> Interpo_5_2:byteenable
	wire  [31:0] mm_interconnect_0_interpo_5_3_s1_writedata;       // mm_interconnect_0:Interpo_5_3_s1_writedata -> Interpo_5_3:writedata
	wire   [5:0] mm_interconnect_0_interpo_5_3_s1_address;         // mm_interconnect_0:Interpo_5_3_s1_address -> Interpo_5_3:address
	wire         mm_interconnect_0_interpo_5_3_s1_chipselect;      // mm_interconnect_0:Interpo_5_3_s1_chipselect -> Interpo_5_3:chipselect
	wire         mm_interconnect_0_interpo_5_3_s1_clken;           // mm_interconnect_0:Interpo_5_3_s1_clken -> Interpo_5_3:clken
	wire         mm_interconnect_0_interpo_5_3_s1_write;           // mm_interconnect_0:Interpo_5_3_s1_write -> Interpo_5_3:write
	wire  [31:0] mm_interconnect_0_interpo_5_3_s1_readdata;        // Interpo_5_3:readdata -> mm_interconnect_0:Interpo_5_3_s1_readdata
	wire   [3:0] mm_interconnect_0_interpo_5_3_s1_byteenable;      // mm_interconnect_0:Interpo_5_3_s1_byteenable -> Interpo_5_3:byteenable
	wire  [31:0] mm_interconnect_0_adapt_fir_mem_s1_writedata;     // mm_interconnect_0:Adapt_FIR_mem_s1_writedata -> Adapt_FIR_mem:writedata
	wire   [8:0] mm_interconnect_0_adapt_fir_mem_s1_address;       // mm_interconnect_0:Adapt_FIR_mem_s1_address -> Adapt_FIR_mem:address
	wire         mm_interconnect_0_adapt_fir_mem_s1_chipselect;    // mm_interconnect_0:Adapt_FIR_mem_s1_chipselect -> Adapt_FIR_mem:chipselect
	wire         mm_interconnect_0_adapt_fir_mem_s1_clken;         // mm_interconnect_0:Adapt_FIR_mem_s1_clken -> Adapt_FIR_mem:clken
	wire         mm_interconnect_0_adapt_fir_mem_s1_write;         // mm_interconnect_0:Adapt_FIR_mem_s1_write -> Adapt_FIR_mem:write
	wire  [31:0] mm_interconnect_0_adapt_fir_mem_s1_readdata;      // Adapt_FIR_mem:readdata -> mm_interconnect_0:Adapt_FIR_mem_s1_readdata
	wire   [3:0] mm_interconnect_0_adapt_fir_mem_s1_byteenable;    // mm_interconnect_0:Adapt_FIR_mem_s1_byteenable -> Adapt_FIR_mem:byteenable
	wire  [31:0] mm_interconnect_0_micfilter_cntl_s1_writedata;    // mm_interconnect_0:micFilter_cntl_s1_writedata -> micFilter_cntl:writedata
	wire   [2:0] mm_interconnect_0_micfilter_cntl_s1_address;      // mm_interconnect_0:micFilter_cntl_s1_address -> micFilter_cntl:address
	wire         mm_interconnect_0_micfilter_cntl_s1_chipselect;   // mm_interconnect_0:micFilter_cntl_s1_chipselect -> micFilter_cntl:chipselect
	wire         mm_interconnect_0_micfilter_cntl_s1_write;        // mm_interconnect_0:micFilter_cntl_s1_write -> micFilter_cntl:write_n
	wire  [31:0] mm_interconnect_0_micfilter_cntl_s1_readdata;     // micFilter_cntl:readdata -> mm_interconnect_0:micFilter_cntl_s1_readdata
	wire  [31:0] mm_interconnect_0_micfilter_rst_s1_writedata;     // mm_interconnect_0:micFilter_rst_s1_writedata -> micFilter_rst:writedata
	wire   [1:0] mm_interconnect_0_micfilter_rst_s1_address;       // mm_interconnect_0:micFilter_rst_s1_address -> micFilter_rst:address
	wire         mm_interconnect_0_micfilter_rst_s1_chipselect;    // mm_interconnect_0:micFilter_rst_s1_chipselect -> micFilter_rst:chipselect
	wire         mm_interconnect_0_micfilter_rst_s1_write;         // mm_interconnect_0:micFilter_rst_s1_write -> micFilter_rst:write_n
	wire  [31:0] mm_interconnect_0_micfilter_rst_s1_readdata;      // micFilter_rst:readdata -> mm_interconnect_0:micFilter_rst_s1_readdata
	wire  [31:0] mm_interconnect_0_micfilter_adjust_s1_writedata;  // mm_interconnect_0:micFilter_adjust_s1_writedata -> micFilter_adjust:writedata
	wire   [1:0] mm_interconnect_0_micfilter_adjust_s1_address;    // mm_interconnect_0:micFilter_adjust_s1_address -> micFilter_adjust:address
	wire         mm_interconnect_0_micfilter_adjust_s1_chipselect; // mm_interconnect_0:micFilter_adjust_s1_chipselect -> micFilter_adjust:chipselect
	wire         mm_interconnect_0_micfilter_adjust_s1_write;      // mm_interconnect_0:micFilter_adjust_s1_write -> micFilter_adjust:write_n
	wire  [31:0] mm_interconnect_0_micfilter_adjust_s1_readdata;   // micFilter_adjust:readdata -> mm_interconnect_0:micFilter_adjust_s1_readdata
	wire  [31:0] mm_interconnect_0_output1_sel_s1_writedata;       // mm_interconnect_0:output1_sel_s1_writedata -> output1_sel:writedata
	wire   [1:0] mm_interconnect_0_output1_sel_s1_address;         // mm_interconnect_0:output1_sel_s1_address -> output1_sel:address
	wire         mm_interconnect_0_output1_sel_s1_chipselect;      // mm_interconnect_0:output1_sel_s1_chipselect -> output1_sel:chipselect
	wire         mm_interconnect_0_output1_sel_s1_write;           // mm_interconnect_0:output1_sel_s1_write -> output1_sel:write_n
	wire  [31:0] mm_interconnect_0_output1_sel_s1_readdata;        // output1_sel:readdata -> mm_interconnect_0:output1_sel_s1_readdata
	wire  [31:0] mm_interconnect_0_output2_sel_s1_writedata;       // mm_interconnect_0:output2_sel_s1_writedata -> output2_sel:writedata
	wire   [1:0] mm_interconnect_0_output2_sel_s1_address;         // mm_interconnect_0:output2_sel_s1_address -> output2_sel:address
	wire         mm_interconnect_0_output2_sel_s1_chipselect;      // mm_interconnect_0:output2_sel_s1_chipselect -> output2_sel:chipselect
	wire         mm_interconnect_0_output2_sel_s1_write;           // mm_interconnect_0:output2_sel_s1_write -> output2_sel:write_n
	wire  [31:0] mm_interconnect_0_output2_sel_s1_readdata;        // output2_sel:readdata -> mm_interconnect_0:output2_sel_s1_readdata
	wire  [31:0] mm_interconnect_0_bypass_sel_s1_writedata;        // mm_interconnect_0:bypass_sel_s1_writedata -> bypass_sel:writedata
	wire   [1:0] mm_interconnect_0_bypass_sel_s1_address;          // mm_interconnect_0:bypass_sel_s1_address -> bypass_sel:address
	wire         mm_interconnect_0_bypass_sel_s1_chipselect;       // mm_interconnect_0:bypass_sel_s1_chipselect -> bypass_sel:chipselect
	wire         mm_interconnect_0_bypass_sel_s1_write;            // mm_interconnect_0:bypass_sel_s1_write -> bypass_sel:write_n
	wire  [31:0] mm_interconnect_0_bypass_sel_s1_readdata;         // bypass_sel:readdata -> mm_interconnect_0:bypass_sel_s1_readdata
	wire  [31:0] mm_interconnect_0_sub_factor_s1_writedata;        // mm_interconnect_0:sub_factor_s1_writedata -> sub_factor:writedata
	wire   [1:0] mm_interconnect_0_sub_factor_s1_address;          // mm_interconnect_0:sub_factor_s1_address -> sub_factor:address
	wire         mm_interconnect_0_sub_factor_s1_chipselect;       // mm_interconnect_0:sub_factor_s1_chipselect -> sub_factor:chipselect
	wire         mm_interconnect_0_sub_factor_s1_write;            // mm_interconnect_0:sub_factor_s1_write -> sub_factor:write_n
	wire  [31:0] mm_interconnect_0_sub_factor_s1_readdata;         // sub_factor:readdata -> mm_interconnect_0:sub_factor_s1_readdata
	wire  [31:0] mm_interconnect_0_delay_lenght_s1_writedata;      // mm_interconnect_0:delay_lenght_s1_writedata -> delay_lenght:writedata
	wire   [1:0] mm_interconnect_0_delay_lenght_s1_address;        // mm_interconnect_0:delay_lenght_s1_address -> delay_lenght:address
	wire         mm_interconnect_0_delay_lenght_s1_chipselect;     // mm_interconnect_0:delay_lenght_s1_chipselect -> delay_lenght:chipselect
	wire         mm_interconnect_0_delay_lenght_s1_write;          // mm_interconnect_0:delay_lenght_s1_write -> delay_lenght:write_n
	wire  [31:0] mm_interconnect_0_delay_lenght_s1_readdata;       // delay_lenght:readdata -> mm_interconnect_0:delay_lenght_s1_readdata
	wire  [31:0] mm_interconnect_0_adapt_pth_s1_writedata;         // mm_interconnect_0:adapt_pTh_s1_writedata -> adapt_pTh:writedata
	wire   [1:0] mm_interconnect_0_adapt_pth_s1_address;           // mm_interconnect_0:adapt_pTh_s1_address -> adapt_pTh:address
	wire         mm_interconnect_0_adapt_pth_s1_chipselect;        // mm_interconnect_0:adapt_pTh_s1_chipselect -> adapt_pTh:chipselect
	wire         mm_interconnect_0_adapt_pth_s1_write;             // mm_interconnect_0:adapt_pTh_s1_write -> adapt_pTh:write_n
	wire  [31:0] mm_interconnect_0_adapt_pth_s1_readdata;          // adapt_pTh:readdata -> mm_interconnect_0:adapt_pTh_s1_readdata
	wire  [31:0] mm_interconnect_0_adapt_weight_s1_writedata;      // mm_interconnect_0:adapt_weight_s1_writedata -> adapt_weight:writedata
	wire   [1:0] mm_interconnect_0_adapt_weight_s1_address;        // mm_interconnect_0:adapt_weight_s1_address -> adapt_weight:address
	wire         mm_interconnect_0_adapt_weight_s1_chipselect;     // mm_interconnect_0:adapt_weight_s1_chipselect -> adapt_weight:chipselect
	wire         mm_interconnect_0_adapt_weight_s1_write;          // mm_interconnect_0:adapt_weight_s1_write -> adapt_weight:write_n
	wire  [31:0] mm_interconnect_0_adapt_weight_s1_readdata;       // adapt_weight:readdata -> mm_interconnect_0:adapt_weight_s1_readdata
	wire  [31:0] mm_interconnect_0_downsamplemult_s1_writedata;    // mm_interconnect_0:DownSampleMult_s1_writedata -> DownSampleMult:writedata
	wire   [1:0] mm_interconnect_0_downsamplemult_s1_address;      // mm_interconnect_0:DownSampleMult_s1_address -> DownSampleMult:address
	wire         mm_interconnect_0_downsamplemult_s1_chipselect;   // mm_interconnect_0:DownSampleMult_s1_chipselect -> DownSampleMult:chipselect
	wire         mm_interconnect_0_downsamplemult_s1_write;        // mm_interconnect_0:DownSampleMult_s1_write -> DownSampleMult:write_n
	wire  [31:0] mm_interconnect_0_downsamplemult_s1_readdata;     // DownSampleMult:readdata -> mm_interconnect_0:DownSampleMult_s1_readdata
	wire  [31:0] mm_interconnect_0_adapt_nth_s1_writedata;         // mm_interconnect_0:adapt_nTh_s1_writedata -> adapt_nTh:writedata
	wire   [1:0] mm_interconnect_0_adapt_nth_s1_address;           // mm_interconnect_0:adapt_nTh_s1_address -> adapt_nTh:address
	wire         mm_interconnect_0_adapt_nth_s1_chipselect;        // mm_interconnect_0:adapt_nTh_s1_chipselect -> adapt_nTh:chipselect
	wire         mm_interconnect_0_adapt_nth_s1_write;             // mm_interconnect_0:adapt_nTh_s1_write -> adapt_nTh:write_n
	wire  [31:0] mm_interconnect_0_adapt_nth_s1_readdata;          // adapt_nTh:readdata -> mm_interconnect_0:adapt_nTh_s1_readdata
	wire         mm_interconnect_0_pcie_ip_txs_waitrequest;        // pcie_ip:txs_waitrequest -> mm_interconnect_0:pcie_ip_txs_waitrequest
	wire   [6:0] mm_interconnect_0_pcie_ip_txs_burstcount;         // mm_interconnect_0:pcie_ip_txs_burstcount -> pcie_ip:txs_burstcount
	wire  [63:0] mm_interconnect_0_pcie_ip_txs_writedata;          // mm_interconnect_0:pcie_ip_txs_writedata -> pcie_ip:txs_writedata
	wire  [30:0] mm_interconnect_0_pcie_ip_txs_address;            // mm_interconnect_0:pcie_ip_txs_address -> pcie_ip:txs_address
	wire         mm_interconnect_0_pcie_ip_txs_chipselect;         // mm_interconnect_0:pcie_ip_txs_chipselect -> pcie_ip:txs_chipselect
	wire         mm_interconnect_0_pcie_ip_txs_write;              // mm_interconnect_0:pcie_ip_txs_write -> pcie_ip:txs_write
	wire         mm_interconnect_0_pcie_ip_txs_read;               // mm_interconnect_0:pcie_ip_txs_read -> pcie_ip:txs_read
	wire  [63:0] mm_interconnect_0_pcie_ip_txs_readdata;           // pcie_ip:txs_readdata -> mm_interconnect_0:pcie_ip_txs_readdata
	wire         mm_interconnect_0_pcie_ip_txs_readdatavalid;      // pcie_ip:txs_readdatavalid -> mm_interconnect_0:pcie_ip_txs_readdatavalid
	wire   [7:0] mm_interconnect_0_pcie_ip_txs_byteenable;         // mm_interconnect_0:pcie_ip_txs_byteenable -> pcie_ip:txs_byteenable
	wire   [6:0] pcie_ip_bar2_burstcount;                          // pcie_ip:bar2_burstcount -> mm_interconnect_1:pcie_ip_bar2_burstcount
	wire         pcie_ip_bar2_waitrequest;                         // mm_interconnect_1:pcie_ip_bar2_waitrequest -> pcie_ip:bar2_waitrequest
	wire  [63:0] pcie_ip_bar2_writedata;                           // pcie_ip:bar2_writedata -> mm_interconnect_1:pcie_ip_bar2_writedata
	wire  [31:0] pcie_ip_bar2_address;                             // pcie_ip:bar2_address -> mm_interconnect_1:pcie_ip_bar2_address
	wire         pcie_ip_bar2_write;                               // pcie_ip:bar2_write -> mm_interconnect_1:pcie_ip_bar2_write
	wire         pcie_ip_bar2_read;                                // pcie_ip:bar2_read -> mm_interconnect_1:pcie_ip_bar2_read
	wire  [63:0] pcie_ip_bar2_readdata;                            // mm_interconnect_1:pcie_ip_bar2_readdata -> pcie_ip:bar2_readdata
	wire   [7:0] pcie_ip_bar2_byteenable;                          // pcie_ip:bar2_byteenable -> mm_interconnect_1:pcie_ip_bar2_byteenable
	wire         pcie_ip_bar2_readdatavalid;                       // mm_interconnect_1:pcie_ip_bar2_readdatavalid -> pcie_ip:bar2_readdatavalid
	wire  [31:0] mm_interconnect_1_sgdma_csr_writedata;            // mm_interconnect_1:sgdma_csr_writedata -> sgdma:csr_writedata
	wire   [3:0] mm_interconnect_1_sgdma_csr_address;              // mm_interconnect_1:sgdma_csr_address -> sgdma:csr_address
	wire         mm_interconnect_1_sgdma_csr_chipselect;           // mm_interconnect_1:sgdma_csr_chipselect -> sgdma:csr_chipselect
	wire         mm_interconnect_1_sgdma_csr_write;                // mm_interconnect_1:sgdma_csr_write -> sgdma:csr_write
	wire         mm_interconnect_1_sgdma_csr_read;                 // mm_interconnect_1:sgdma_csr_read -> sgdma:csr_read
	wire  [31:0] mm_interconnect_1_sgdma_csr_readdata;             // sgdma:csr_readdata -> mm_interconnect_1:sgdma_csr_readdata
	wire         mm_interconnect_1_pcie_ip_cra_waitrequest;        // pcie_ip:cra_waitrequest -> mm_interconnect_1:pcie_ip_cra_waitrequest
	wire  [31:0] mm_interconnect_1_pcie_ip_cra_writedata;          // mm_interconnect_1:pcie_ip_cra_writedata -> pcie_ip:cra_writedata
	wire  [11:0] mm_interconnect_1_pcie_ip_cra_address;            // mm_interconnect_1:pcie_ip_cra_address -> pcie_ip:cra_address
	wire         mm_interconnect_1_pcie_ip_cra_chipselect;         // mm_interconnect_1:pcie_ip_cra_chipselect -> pcie_ip:cra_chipselect
	wire         mm_interconnect_1_pcie_ip_cra_write;              // mm_interconnect_1:pcie_ip_cra_write -> pcie_ip:cra_write
	wire         mm_interconnect_1_pcie_ip_cra_read;               // mm_interconnect_1:pcie_ip_cra_read -> pcie_ip:cra_read
	wire  [31:0] mm_interconnect_1_pcie_ip_cra_readdata;           // pcie_ip:cra_readdata -> mm_interconnect_1:pcie_ip_cra_readdata
	wire   [3:0] mm_interconnect_1_pcie_ip_cra_byteenable;         // mm_interconnect_1:pcie_ip_cra_byteenable -> pcie_ip:cra_byteenable
	wire         irq_mapper_receiver0_irq;                         // sgdma:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                         // fifo_memory:wrclk_control_slave_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                         // button:irq -> irq_mapper:receiver2_irq
	wire  [15:0] pcie_ip_rxm_irq_irq;                              // irq_mapper:sender_irq -> pcie_ip:rxm_irq_irq
	wire         rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [Adapt_FIR_mem:reset, DownSampleMult:reset_n, Interpo_4_0:reset, Interpo_5_0:reset, Interpo_5_1:reset, Interpo_5_2:reset, Interpo_5_3:reset, adapt_nTh:reset_n, adapt_pTh:reset_n, adapt_weight:reset_n, button:reset_n, bypass_sel:reset_n, delay_lenght:reset_n, fifo_memory:reset_n, fir_memory:reset, led:reset_n, micFilter_adjust:reset_n, micFilter_cntl:reset_n, micFilter_rst:reset_n, mm_interconnect_0:sgdma_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sgdma_reset_reset_bridge_in_reset_reset, output1_sel:reset_n, output2_sel:reset_n, rst_translator:in_reset, sgdma:system_reset_n, sub_factor:reset_n]
	wire         rst_controller_reset_out_reset_req;               // rst_controller:reset_req -> [Adapt_FIR_mem:reset_req, Interpo_4_0:reset_req, Interpo_5_0:reset_req, Interpo_5_1:reset_req, Interpo_5_2:reset_req, Interpo_5_3:reset_req, fir_memory:reset_req, rst_translator:reset_req_in]
	wire         pcie_ip_pcie_core_reset_reset;                    // pcie_ip:pcie_core_reset_reset_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;               // rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pcie_ip_bar2_translator_reset_reset_bridge_in_reset_reset]

	de2i_150_qsys_pcie_ip #(
		.p_pcie_hip_type                     ("2"),
		.lane_mask                           (8'b11111110),
		.max_link_width                      (1),
		.millisecond_cycle_count             ("125000"),
		.enable_gen2_core                    ("false"),
		.gen2_lane_rate_mode                 ("false"),
		.no_soft_reset                       ("false"),
		.core_clk_divider                    (2),
		.enable_ch0_pclk_out                 ("true"),
		.core_clk_source                     ("pclk"),
		.CB_P2A_AVALON_ADDR_B0               (0),
		.bar0_size_mask                      (19),
		.bar0_io_space                       ("false"),
		.bar0_64bit_mem_space                ("true"),
		.bar0_prefetchable                   ("true"),
		.CB_P2A_AVALON_ADDR_B1               (0),
		.bar1_size_mask                      (0),
		.bar1_io_space                       ("false"),
		.bar1_64bit_mem_space                ("true"),
		.bar1_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B2               (0),
		.bar2_size_mask                      (15),
		.bar2_io_space                       ("false"),
		.bar2_64bit_mem_space                ("false"),
		.bar2_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B3               (0),
		.bar3_size_mask                      (0),
		.bar3_io_space                       ("false"),
		.bar3_64bit_mem_space                ("false"),
		.bar3_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B4               (0),
		.bar4_size_mask                      (0),
		.bar4_io_space                       ("false"),
		.bar4_64bit_mem_space                ("false"),
		.bar4_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B5               (0),
		.bar5_size_mask                      (0),
		.bar5_io_space                       ("false"),
		.bar5_64bit_mem_space                ("false"),
		.bar5_prefetchable                   ("false"),
		.vendor_id                           (4466),
		.device_id                           (57345),
		.revision_id                         (1),
		.class_code                          (0),
		.subsystem_vendor_id                 (4466),
		.subsystem_device_id                 (4),
		.port_link_number                    (1),
		.msi_function_count                  (0),
		.enable_msi_64bit_addressing         ("true"),
		.enable_function_msix_support        ("false"),
		.eie_before_nfts_count               (4),
		.enable_completion_timeout_disable   ("false"),
		.completion_timeout                  ("NONE"),
		.enable_adapter_half_rate_mode       ("false"),
		.msix_pba_bir                        (0),
		.msix_pba_offset                     (0),
		.msix_table_bir                      (0),
		.msix_table_offset                   (0),
		.msix_table_size                     (0),
		.use_crc_forwarding                  ("false"),
		.surprise_down_error_support         ("false"),
		.dll_active_report_support           ("false"),
		.bar_io_window_size                  ("32BIT"),
		.bar_prefetchable                    (32),
		.hot_plug_support                    (7'b0000000),
		.no_command_completed                ("true"),
		.slot_power_limit                    (0),
		.slot_power_scale                    (0),
		.slot_number                         (0),
		.enable_slot_register                ("false"),
		.advanced_errors                     ("false"),
		.enable_ecrc_check                   ("false"),
		.enable_ecrc_gen                     ("false"),
		.max_payload_size                    (0),
		.retry_buffer_last_active_address    (255),
		.credit_buffer_allocation_aux        ("ABSOLUTE"),
		.vc0_rx_flow_ctrl_posted_header      (28),
		.vc0_rx_flow_ctrl_posted_data        (198),
		.vc0_rx_flow_ctrl_nonposted_header   (30),
		.vc0_rx_flow_ctrl_nonposted_data     (0),
		.vc0_rx_flow_ctrl_compl_header       (48),
		.vc0_rx_flow_ctrl_compl_data         (256),
		.RX_BUF                              (9),
		.RH_NUM                              (7),
		.G_TAG_NUM0                          (32),
		.endpoint_l0_latency                 (0),
		.endpoint_l1_latency                 (0),
		.enable_l1_aspm                      ("false"),
		.l01_entry_latency                   (31),
		.diffclock_nfts_count                (255),
		.sameclock_nfts_count                (255),
		.l1_exit_latency_sameclock           (7),
		.l1_exit_latency_diffclock           (7),
		.l0_exit_latency_sameclock           (7),
		.l0_exit_latency_diffclock           (7),
		.gen2_diffclock_nfts_count           (255),
		.gen2_sameclock_nfts_count           (255),
		.CG_COMMON_CLOCK_MODE                (1),
		.CB_PCIE_MODE                        (0),
		.AST_LITE                            (0),
		.CB_PCIE_RX_LITE                     (0),
		.CG_RXM_IRQ_NUM                      (16),
		.CG_AVALON_S_ADDR_WIDTH              (20),
		.bypass_tl                           ("false"),
		.CG_IMPL_CRA_AV_SLAVE_PORT           (1),
		.CG_NO_CPL_REORDERING                (0),
		.CG_ENABLE_A2P_INTERRUPT             (0),
		.p_user_msi_enable                   (0),
		.CG_IRQ_BIT_ENA                      (65535),
		.CB_A2P_ADDR_MAP_IS_FIXED            (1),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES         (1),
		.CB_A2P_ADDR_MAP_PASS_THRU_BITS      (31),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_LOW  (32'b00000000000000000000000000000000),
		.RXM_DATA_WIDTH                      (64),
		.RXM_BEN_WIDTH                       (8),
		.TL_SELECTION                        (1),
		.pcie_mode                           ("SHARED_MODE"),
		.single_rx_detect                    (1),
		.enable_coreclk_out_half_rate        ("false"),
		.low_priority_vc                     (0),
		.link_width                          (1),
		.cyclone4                            (1)
	) pcie_ip (
		.pcie_core_clk_clk                  (pcie_ip_pcie_core_clk_clk),                   //      pcie_core_clk.clk
		.pcie_core_reset_reset_n            (pcie_ip_pcie_core_reset_reset),               //    pcie_core_reset.reset_n
		.cal_blk_clk_clk                    (clk_clk),                                     //        cal_blk_clk.clk
		.txs_address                        (mm_interconnect_0_pcie_ip_txs_address),       //                txs.address
		.txs_chipselect                     (mm_interconnect_0_pcie_ip_txs_chipselect),    //                   .chipselect
		.txs_byteenable                     (mm_interconnect_0_pcie_ip_txs_byteenable),    //                   .byteenable
		.txs_readdata                       (mm_interconnect_0_pcie_ip_txs_readdata),      //                   .readdata
		.txs_writedata                      (mm_interconnect_0_pcie_ip_txs_writedata),     //                   .writedata
		.txs_read                           (mm_interconnect_0_pcie_ip_txs_read),          //                   .read
		.txs_write                          (mm_interconnect_0_pcie_ip_txs_write),         //                   .write
		.txs_burstcount                     (mm_interconnect_0_pcie_ip_txs_burstcount),    //                   .burstcount
		.txs_readdatavalid                  (mm_interconnect_0_pcie_ip_txs_readdatavalid), //                   .readdatavalid
		.txs_waitrequest                    (mm_interconnect_0_pcie_ip_txs_waitrequest),   //                   .waitrequest
		.refclk_export                      (pcie_ip_refclk_export),                       //             refclk.export
		.test_in_test_in                    (pcie_ip_test_in_test_in),                     //            test_in.test_in
		.pcie_rstn_export                   (pcie_ip_pcie_rstn_export),                    //          pcie_rstn.export
		.clocks_sim_clk250_export           (pcie_ip_clocks_sim_clk250_export),            //         clocks_sim.clk250_export
		.clocks_sim_clk500_export           (pcie_ip_clocks_sim_clk500_export),            //                   .clk500_export
		.clocks_sim_clk125_export           (pcie_ip_clocks_sim_clk125_export),            //                   .clk125_export
		.reconfig_busy_busy_altgxb_reconfig (pcie_ip_reconfig_busy_busy_altgxb_reconfig),  //      reconfig_busy.busy_altgxb_reconfig
		.pipe_ext_pipe_mode                 (pcie_ip_pipe_ext_pipe_mode),                  //           pipe_ext.pipe_mode
		.pipe_ext_phystatus_ext             (pcie_ip_pipe_ext_phystatus_ext),              //                   .phystatus_ext
		.pipe_ext_rate_ext                  (pcie_ip_pipe_ext_rate_ext),                   //                   .rate_ext
		.pipe_ext_powerdown_ext             (pcie_ip_pipe_ext_powerdown_ext),              //                   .powerdown_ext
		.pipe_ext_txdetectrx_ext            (pcie_ip_pipe_ext_txdetectrx_ext),             //                   .txdetectrx_ext
		.pipe_ext_rxelecidle0_ext           (pcie_ip_pipe_ext_rxelecidle0_ext),            //                   .rxelecidle0_ext
		.pipe_ext_rxdata0_ext               (pcie_ip_pipe_ext_rxdata0_ext),                //                   .rxdata0_ext
		.pipe_ext_rxstatus0_ext             (pcie_ip_pipe_ext_rxstatus0_ext),              //                   .rxstatus0_ext
		.pipe_ext_rxvalid0_ext              (pcie_ip_pipe_ext_rxvalid0_ext),               //                   .rxvalid0_ext
		.pipe_ext_rxdatak0_ext              (pcie_ip_pipe_ext_rxdatak0_ext),               //                   .rxdatak0_ext
		.pipe_ext_txdata0_ext               (pcie_ip_pipe_ext_txdata0_ext),                //                   .txdata0_ext
		.pipe_ext_txdatak0_ext              (pcie_ip_pipe_ext_txdatak0_ext),               //                   .txdatak0_ext
		.pipe_ext_rxpolarity0_ext           (pcie_ip_pipe_ext_rxpolarity0_ext),            //                   .rxpolarity0_ext
		.pipe_ext_txcompl0_ext              (pcie_ip_pipe_ext_txcompl0_ext),               //                   .txcompl0_ext
		.pipe_ext_txelecidle0_ext           (pcie_ip_pipe_ext_txelecidle0_ext),            //                   .txelecidle0_ext
		.powerdown_pll_powerdown            (),                                            //          powerdown.pll_powerdown
		.powerdown_gxb_powerdown            (),                                            //                   .gxb_powerdown
		.bar1_0_address                     (pcie_ip_bar1_0_address),                      //             bar1_0.address
		.bar1_0_read                        (pcie_ip_bar1_0_read),                         //                   .read
		.bar1_0_waitrequest                 (pcie_ip_bar1_0_waitrequest),                  //                   .waitrequest
		.bar1_0_write                       (pcie_ip_bar1_0_write),                        //                   .write
		.bar1_0_readdatavalid               (pcie_ip_bar1_0_readdatavalid),                //                   .readdatavalid
		.bar1_0_readdata                    (pcie_ip_bar1_0_readdata),                     //                   .readdata
		.bar1_0_writedata                   (pcie_ip_bar1_0_writedata),                    //                   .writedata
		.bar1_0_burstcount                  (pcie_ip_bar1_0_burstcount),                   //                   .burstcount
		.bar1_0_byteenable                  (pcie_ip_bar1_0_byteenable),                   //                   .byteenable
		.bar2_address                       (pcie_ip_bar2_address),                        //               bar2.address
		.bar2_read                          (pcie_ip_bar2_read),                           //                   .read
		.bar2_waitrequest                   (pcie_ip_bar2_waitrequest),                    //                   .waitrequest
		.bar2_write                         (pcie_ip_bar2_write),                          //                   .write
		.bar2_readdatavalid                 (pcie_ip_bar2_readdatavalid),                  //                   .readdatavalid
		.bar2_readdata                      (pcie_ip_bar2_readdata),                       //                   .readdata
		.bar2_writedata                     (pcie_ip_bar2_writedata),                      //                   .writedata
		.bar2_burstcount                    (pcie_ip_bar2_burstcount),                     //                   .burstcount
		.bar2_byteenable                    (pcie_ip_bar2_byteenable),                     //                   .byteenable
		.cra_chipselect                     (mm_interconnect_1_pcie_ip_cra_chipselect),    //                cra.chipselect
		.cra_address                        (mm_interconnect_1_pcie_ip_cra_address),       //                   .address
		.cra_byteenable                     (mm_interconnect_1_pcie_ip_cra_byteenable),    //                   .byteenable
		.cra_read                           (mm_interconnect_1_pcie_ip_cra_read),          //                   .read
		.cra_readdata                       (mm_interconnect_1_pcie_ip_cra_readdata),      //                   .readdata
		.cra_write                          (mm_interconnect_1_pcie_ip_cra_write),         //                   .write
		.cra_writedata                      (mm_interconnect_1_pcie_ip_cra_writedata),     //                   .writedata
		.cra_waitrequest                    (mm_interconnect_1_pcie_ip_cra_waitrequest),   //                   .waitrequest
		.cra_irq_irq                        (),                                            //            cra_irq.irq
		.rxm_irq_irq                        (pcie_ip_rxm_irq_irq),                         //            rxm_irq.irq
		.rx_in_rx_datain_0                  (pcie_ip_rx_in_rx_datain_0),                   //              rx_in.rx_datain_0
		.tx_out_tx_dataout_0                (pcie_ip_tx_out_tx_dataout_0),                 //             tx_out.tx_dataout_0
		.reconfig_togxb_data                (pcie_ip_reconfig_togxb_data),                 //     reconfig_togxb.data
		.reconfig_gxbclk_clk                (clk_clk),                                     //    reconfig_gxbclk.clk
		.reconfig_fromgxb_0_data            (pcie_ip_reconfig_fromgxb_0_data),             // reconfig_fromgxb_0.data
		.fixedclk_clk                       (pcie_ip_pcie_core_clk_clk)                    //           fixedclk.clk
	);

	de2i_150_qsys_sgdma sgdma (
		.clk                           (pcie_ip_pcie_core_clk_clk),              //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),        //            reset.reset_n
		.csr_chipselect                (mm_interconnect_1_sgdma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_1_sgdma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_1_sgdma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_1_sgdma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_1_sgdma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_1_sgdma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),               //          csr_irq.irq
		.m_read_readdata               (sgdma_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_m_read_read),                      //                 .read
		.m_write_waitrequest           (sgdma_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_m_write_byteenable)                //                 .byteenable
	);

	de2i_150_qsys_fir_memory fir_memory (
		.clk         (pcie_ip_pcie_core_clk_clk),                  //   clk1.clk
		.address     (mm_interconnect_0_fir_memory_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_fir_memory_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_fir_memory_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_fir_memory_s1_write),      //       .write
		.readdata    (mm_interconnect_0_fir_memory_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_fir_memory_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_fir_memory_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),         //       .reset_req
		.address2    (fir_memory_s2_address),                      //     s2.address
		.chipselect2 (fir_memory_s2_chipselect),                   //       .chipselect
		.clken2      (fir_memory_s2_clken),                        //       .clken
		.write2      (fir_memory_s2_write),                        //       .write
		.readdata2   (fir_memory_s2_readdata),                     //       .readdata
		.writedata2  (fir_memory_s2_writedata),                    //       .writedata
		.byteenable2 (fir_memory_s2_byteenable),                   //       .byteenable
		.clk2        (fir_memory_clk2_clk),                        //   clk2.clk
		.reset2      (fir_memory_reset2_reset),                    // reset2.reset
		.reset_req2  (fir_memory_reset2_reset_req)                 //       .reset_req
	);

	de2i_150_qsys_led led (
		.clk        (pcie_ip_pcie_core_clk_clk),           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	de2i_150_qsys_button button (
		.clk        (pcie_ip_pcie_core_clk_clk),              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_button_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_s1_readdata),   //                    .readdata
		.in_port    (button_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                //                 irq.irq
	);

	de2i_150_qsys_fifo_memory fifo_memory (
		.wrclock                          (pcie_ip_pcie_core_clk_clk),                      //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),                // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_memory_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_memory_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_memory_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_memory_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_memory_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_memory_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_memory_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_memory_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_memory_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_memory_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_memory_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver1_irq)                        //   in_irq.irq
	);

	de2i_150_qsys_Interpo_4_0 interpo_4_0 (
		.clk         (pcie_ip_pcie_core_clk_clk),                   //   clk1.clk
		.address     (mm_interconnect_0_interpo_4_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_interpo_4_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_interpo_4_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_interpo_4_0_s1_write),      //       .write
		.readdata    (mm_interconnect_0_interpo_4_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_interpo_4_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_interpo_4_0_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.address2    (interpo_4_0_s2_address),                      //     s2.address
		.chipselect2 (interpo_4_0_s2_chipselect),                   //       .chipselect
		.clken2      (interpo_4_0_s2_clken),                        //       .clken
		.write2      (interpo_4_0_s2_write),                        //       .write
		.readdata2   (interpo_4_0_s2_readdata),                     //       .readdata
		.writedata2  (interpo_4_0_s2_writedata),                    //       .writedata
		.byteenable2 (interpo_4_0_s2_byteenable),                   //       .byteenable
		.clk2        (interpo_4_0_clk2_clk),                        //   clk2.clk
		.reset2      (interpo_4_0_reset2_reset),                    // reset2.reset
		.reset_req2  (interpo_4_0_reset2_reset_req)                 //       .reset_req
	);

	de2i_150_qsys_Interpo_5_0 interpo_5_0 (
		.clk         (pcie_ip_pcie_core_clk_clk),                   //   clk1.clk
		.address     (mm_interconnect_0_interpo_5_0_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_interpo_5_0_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_interpo_5_0_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_interpo_5_0_s1_write),      //       .write
		.readdata    (mm_interconnect_0_interpo_5_0_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_interpo_5_0_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_interpo_5_0_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.address2    (interpo_5_0_s2_address),                      //     s2.address
		.chipselect2 (interpo_5_0_s2_chipselect),                   //       .chipselect
		.clken2      (interpo_5_0_s2_clken),                        //       .clken
		.write2      (interpo_5_0_s2_write),                        //       .write
		.readdata2   (interpo_5_0_s2_readdata),                     //       .readdata
		.writedata2  (interpo_5_0_s2_writedata),                    //       .writedata
		.byteenable2 (interpo_5_0_s2_byteenable),                   //       .byteenable
		.clk2        (interpo_5_0_clk2_clk),                        //   clk2.clk
		.reset2      (interpo_5_0_reset2_reset),                    // reset2.reset
		.reset_req2  (interpo_5_0_reset2_reset_req)                 //       .reset_req
	);

	de2i_150_qsys_Interpo_5_1 interpo_5_1 (
		.clk         (pcie_ip_pcie_core_clk_clk),                   //   clk1.clk
		.address     (mm_interconnect_0_interpo_5_1_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_interpo_5_1_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_interpo_5_1_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_interpo_5_1_s1_write),      //       .write
		.readdata    (mm_interconnect_0_interpo_5_1_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_interpo_5_1_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_interpo_5_1_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.address2    (interpo_5_1_s2_address),                      //     s2.address
		.chipselect2 (interpo_5_1_s2_chipselect),                   //       .chipselect
		.clken2      (interpo_5_1_s2_clken),                        //       .clken
		.write2      (interpo_5_1_s2_write),                        //       .write
		.readdata2   (interpo_5_1_s2_readdata),                     //       .readdata
		.writedata2  (interpo_5_1_s2_writedata),                    //       .writedata
		.byteenable2 (interpo_5_1_s2_byteenable),                   //       .byteenable
		.clk2        (interpo_5_1_clk2_clk),                        //   clk2.clk
		.reset2      (interpo_5_1_reset2_reset),                    // reset2.reset
		.reset_req2  (interpo_5_1_reset2_reset_req)                 //       .reset_req
	);

	de2i_150_qsys_Interpo_5_2 interpo_5_2 (
		.clk         (pcie_ip_pcie_core_clk_clk),                   //   clk1.clk
		.address     (mm_interconnect_0_interpo_5_2_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_interpo_5_2_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_interpo_5_2_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_interpo_5_2_s1_write),      //       .write
		.readdata    (mm_interconnect_0_interpo_5_2_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_interpo_5_2_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_interpo_5_2_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.address2    (interpo_5_2_s2_address),                      //     s2.address
		.chipselect2 (interpo_5_2_s2_chipselect),                   //       .chipselect
		.clken2      (interpo_5_2_s2_clken),                        //       .clken
		.write2      (interpo_5_2_s2_write),                        //       .write
		.readdata2   (interpo_5_2_s2_readdata),                     //       .readdata
		.writedata2  (interpo_5_2_s2_writedata),                    //       .writedata
		.byteenable2 (interpo_5_2_s2_byteenable),                   //       .byteenable
		.clk2        (interpo_5_2_clk2_clk),                        //   clk2.clk
		.reset2      (interpo_5_2_reset2_reset),                    // reset2.reset
		.reset_req2  (interpo_5_2_reset2_reset_req)                 //       .reset_req
	);

	de2i_150_qsys_Interpo_5_3 interpo_5_3 (
		.clk         (pcie_ip_pcie_core_clk_clk),                   //   clk1.clk
		.address     (mm_interconnect_0_interpo_5_3_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_interpo_5_3_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_interpo_5_3_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_interpo_5_3_s1_write),      //       .write
		.readdata    (mm_interconnect_0_interpo_5_3_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_interpo_5_3_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_interpo_5_3_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.address2    (interpo_5_3_s2_address),                      //     s2.address
		.chipselect2 (interpo_5_3_s2_chipselect),                   //       .chipselect
		.clken2      (interpo_5_3_s2_clken),                        //       .clken
		.write2      (interpo_5_3_s2_write),                        //       .write
		.readdata2   (interpo_5_3_s2_readdata),                     //       .readdata
		.writedata2  (interpo_5_3_s2_writedata),                    //       .writedata
		.byteenable2 (interpo_5_3_s2_byteenable),                   //       .byteenable
		.clk2        (interpo_5_3_clk2_clk),                        //   clk2.clk
		.reset2      (interpo_5_3_reset2_reset),                    // reset2.reset
		.reset_req2  (interpo_5_3_reset2_reset_req)                 //       .reset_req
	);

	de2i_150_qsys_Adapt_FIR_mem adapt_fir_mem (
		.clk         (pcie_ip_pcie_core_clk_clk),                     //   clk1.clk
		.address     (mm_interconnect_0_adapt_fir_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_adapt_fir_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_adapt_fir_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_adapt_fir_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_0_adapt_fir_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_adapt_fir_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_adapt_fir_mem_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),            //       .reset_req
		.address2    (adapt_fir_mem_s2_address),                      //     s2.address
		.chipselect2 (adapt_fir_mem_s2_chipselect),                   //       .chipselect
		.clken2      (adapt_fir_mem_s2_clken),                        //       .clken
		.write2      (adapt_fir_mem_s2_write),                        //       .write
		.readdata2   (adapt_fir_mem_s2_readdata),                     //       .readdata
		.writedata2  (adapt_fir_mem_s2_writedata),                    //       .writedata
		.byteenable2 (adapt_fir_mem_s2_byteenable),                   //       .byteenable
		.clk2        (adapt_fir_mem_clk2_clk),                        //   clk2.clk
		.reset2      (adapt_fir_mem_reset2_reset),                    // reset2.reset
		.reset_req2  (adapt_fir_mem_reset2_reset_req)                 //       .reset_req
	);

	de2i_150_qsys_micFilter_cntl micfilter_cntl (
		.clk        (pcie_ip_pcie_core_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_micfilter_cntl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_micfilter_cntl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_micfilter_cntl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_micfilter_cntl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_micfilter_cntl_s1_readdata),   //                    .readdata
		.out_port   (micfilter_cntl_export)                           // external_connection.export
	);

	de2i_150_qsys_micFilter_rst micfilter_rst (
		.clk        (pcie_ip_pcie_core_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_micfilter_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_micfilter_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_micfilter_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_micfilter_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_micfilter_rst_s1_readdata),   //                    .readdata
		.out_port   (micfilter_rst_export)                           // external_connection.export
	);

	de2i_150_qsys_micFilter_rst micfilter_adjust (
		.clk        (pcie_ip_pcie_core_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_micfilter_adjust_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_micfilter_adjust_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_micfilter_adjust_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_micfilter_adjust_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_micfilter_adjust_s1_readdata),   //                    .readdata
		.out_port   (micfilter_adjust_export)                           // external_connection.export
	);

	de2i_150_qsys_led output1_sel (
		.clk        (pcie_ip_pcie_core_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_output1_sel_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_output1_sel_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_output1_sel_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_output1_sel_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_output1_sel_s1_readdata),   //                    .readdata
		.out_port   (output1_sel_export)                           // external_connection.export
	);

	de2i_150_qsys_led output2_sel (
		.clk        (pcie_ip_pcie_core_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_output2_sel_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_output2_sel_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_output2_sel_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_output2_sel_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_output2_sel_s1_readdata),   //                    .readdata
		.out_port   (output2_sel_export)                           // external_connection.export
	);

	de2i_150_qsys_bypass_sel bypass_sel (
		.clk        (pcie_ip_pcie_core_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_bypass_sel_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bypass_sel_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bypass_sel_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bypass_sel_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bypass_sel_s1_readdata),   //                    .readdata
		.out_port   (bypass_sel_export)                           // external_connection.export
	);

	de2i_150_qsys_sub_factor sub_factor (
		.clk        (pcie_ip_pcie_core_clk_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_sub_factor_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sub_factor_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sub_factor_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sub_factor_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sub_factor_s1_readdata),   //                    .readdata
		.out_port   (sub_factor_export)                           // external_connection.export
	);

	de2i_150_qsys_delay_lenght delay_lenght (
		.clk        (pcie_ip_pcie_core_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_delay_lenght_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_delay_lenght_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_delay_lenght_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_delay_lenght_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_delay_lenght_s1_readdata),   //                    .readdata
		.out_port   (delay_lenght_export)                           // external_connection.export
	);

	de2i_150_qsys_DownSampleMult downsamplemult (
		.clk        (pcie_ip_pcie_core_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_downsamplemult_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_downsamplemult_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_downsamplemult_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_downsamplemult_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_downsamplemult_s1_readdata),   //                    .readdata
		.out_port   (downsamplemult_export)                           // external_connection.export
	);

	de2i_150_qsys_DownSampleMult adapt_weight (
		.clk        (pcie_ip_pcie_core_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_adapt_weight_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_adapt_weight_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_adapt_weight_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_adapt_weight_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_adapt_weight_s1_readdata),   //                    .readdata
		.out_port   (adapt_weight_export)                           // external_connection.export
	);

	de2i_150_qsys_sub_factor adapt_pth (
		.clk        (pcie_ip_pcie_core_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_adapt_pth_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_adapt_pth_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_adapt_pth_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_adapt_pth_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_adapt_pth_s1_readdata),   //                    .readdata
		.out_port   (adapt_pth_export)                           // external_connection.export
	);

	de2i_150_qsys_sub_factor adapt_nth (
		.clk        (pcie_ip_pcie_core_clk_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_adapt_nth_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_adapt_nth_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_adapt_nth_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_adapt_nth_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_adapt_nth_s1_readdata),   //                    .readdata
		.out_port   (adapt_nth_export)                           // external_connection.export
	);

	de2i_150_qsys_mm_interconnect_0 mm_interconnect_0 (
		.pcie_ip_pcie_core_clk_clk                                   (pcie_ip_pcie_core_clk_clk),                        //                                 pcie_ip_pcie_core_clk.clk
		.pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),               // pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset.reset
		.sgdma_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                   //                     sgdma_reset_reset_bridge_in_reset.reset
		.pcie_ip_bar1_0_address                                      (pcie_ip_bar1_0_address),                           //                                        pcie_ip_bar1_0.address
		.pcie_ip_bar1_0_waitrequest                                  (pcie_ip_bar1_0_waitrequest),                       //                                                      .waitrequest
		.pcie_ip_bar1_0_burstcount                                   (pcie_ip_bar1_0_burstcount),                        //                                                      .burstcount
		.pcie_ip_bar1_0_byteenable                                   (pcie_ip_bar1_0_byteenable),                        //                                                      .byteenable
		.pcie_ip_bar1_0_read                                         (pcie_ip_bar1_0_read),                              //                                                      .read
		.pcie_ip_bar1_0_readdata                                     (pcie_ip_bar1_0_readdata),                          //                                                      .readdata
		.pcie_ip_bar1_0_readdatavalid                                (pcie_ip_bar1_0_readdatavalid),                     //                                                      .readdatavalid
		.pcie_ip_bar1_0_write                                        (pcie_ip_bar1_0_write),                             //                                                      .write
		.pcie_ip_bar1_0_writedata                                    (pcie_ip_bar1_0_writedata),                         //                                                      .writedata
		.sgdma_descriptor_read_address                               (sgdma_descriptor_read_address),                    //                                 sgdma_descriptor_read.address
		.sgdma_descriptor_read_waitrequest                           (sgdma_descriptor_read_waitrequest),                //                                                      .waitrequest
		.sgdma_descriptor_read_read                                  (sgdma_descriptor_read_read),                       //                                                      .read
		.sgdma_descriptor_read_readdata                              (sgdma_descriptor_read_readdata),                   //                                                      .readdata
		.sgdma_descriptor_read_readdatavalid                         (sgdma_descriptor_read_readdatavalid),              //                                                      .readdatavalid
		.sgdma_descriptor_write_address                              (sgdma_descriptor_write_address),                   //                                sgdma_descriptor_write.address
		.sgdma_descriptor_write_waitrequest                          (sgdma_descriptor_write_waitrequest),               //                                                      .waitrequest
		.sgdma_descriptor_write_write                                (sgdma_descriptor_write_write),                     //                                                      .write
		.sgdma_descriptor_write_writedata                            (sgdma_descriptor_write_writedata),                 //                                                      .writedata
		.sgdma_m_read_address                                        (sgdma_m_read_address),                             //                                          sgdma_m_read.address
		.sgdma_m_read_waitrequest                                    (sgdma_m_read_waitrequest),                         //                                                      .waitrequest
		.sgdma_m_read_read                                           (sgdma_m_read_read),                                //                                                      .read
		.sgdma_m_read_readdata                                       (sgdma_m_read_readdata),                            //                                                      .readdata
		.sgdma_m_read_readdatavalid                                  (sgdma_m_read_readdatavalid),                       //                                                      .readdatavalid
		.sgdma_m_write_address                                       (sgdma_m_write_address),                            //                                         sgdma_m_write.address
		.sgdma_m_write_waitrequest                                   (sgdma_m_write_waitrequest),                        //                                                      .waitrequest
		.sgdma_m_write_byteenable                                    (sgdma_m_write_byteenable),                         //                                                      .byteenable
		.sgdma_m_write_write                                         (sgdma_m_write_write),                              //                                                      .write
		.sgdma_m_write_writedata                                     (sgdma_m_write_writedata),                          //                                                      .writedata
		.Adapt_FIR_mem_s1_address                                    (mm_interconnect_0_adapt_fir_mem_s1_address),       //                                      Adapt_FIR_mem_s1.address
		.Adapt_FIR_mem_s1_write                                      (mm_interconnect_0_adapt_fir_mem_s1_write),         //                                                      .write
		.Adapt_FIR_mem_s1_readdata                                   (mm_interconnect_0_adapt_fir_mem_s1_readdata),      //                                                      .readdata
		.Adapt_FIR_mem_s1_writedata                                  (mm_interconnect_0_adapt_fir_mem_s1_writedata),     //                                                      .writedata
		.Adapt_FIR_mem_s1_byteenable                                 (mm_interconnect_0_adapt_fir_mem_s1_byteenable),    //                                                      .byteenable
		.Adapt_FIR_mem_s1_chipselect                                 (mm_interconnect_0_adapt_fir_mem_s1_chipselect),    //                                                      .chipselect
		.Adapt_FIR_mem_s1_clken                                      (mm_interconnect_0_adapt_fir_mem_s1_clken),         //                                                      .clken
		.adapt_nTh_s1_address                                        (mm_interconnect_0_adapt_nth_s1_address),           //                                          adapt_nTh_s1.address
		.adapt_nTh_s1_write                                          (mm_interconnect_0_adapt_nth_s1_write),             //                                                      .write
		.adapt_nTh_s1_readdata                                       (mm_interconnect_0_adapt_nth_s1_readdata),          //                                                      .readdata
		.adapt_nTh_s1_writedata                                      (mm_interconnect_0_adapt_nth_s1_writedata),         //                                                      .writedata
		.adapt_nTh_s1_chipselect                                     (mm_interconnect_0_adapt_nth_s1_chipselect),        //                                                      .chipselect
		.adapt_pTh_s1_address                                        (mm_interconnect_0_adapt_pth_s1_address),           //                                          adapt_pTh_s1.address
		.adapt_pTh_s1_write                                          (mm_interconnect_0_adapt_pth_s1_write),             //                                                      .write
		.adapt_pTh_s1_readdata                                       (mm_interconnect_0_adapt_pth_s1_readdata),          //                                                      .readdata
		.adapt_pTh_s1_writedata                                      (mm_interconnect_0_adapt_pth_s1_writedata),         //                                                      .writedata
		.adapt_pTh_s1_chipselect                                     (mm_interconnect_0_adapt_pth_s1_chipselect),        //                                                      .chipselect
		.adapt_weight_s1_address                                     (mm_interconnect_0_adapt_weight_s1_address),        //                                       adapt_weight_s1.address
		.adapt_weight_s1_write                                       (mm_interconnect_0_adapt_weight_s1_write),          //                                                      .write
		.adapt_weight_s1_readdata                                    (mm_interconnect_0_adapt_weight_s1_readdata),       //                                                      .readdata
		.adapt_weight_s1_writedata                                   (mm_interconnect_0_adapt_weight_s1_writedata),      //                                                      .writedata
		.adapt_weight_s1_chipselect                                  (mm_interconnect_0_adapt_weight_s1_chipselect),     //                                                      .chipselect
		.button_s1_address                                           (mm_interconnect_0_button_s1_address),              //                                             button_s1.address
		.button_s1_write                                             (mm_interconnect_0_button_s1_write),                //                                                      .write
		.button_s1_readdata                                          (mm_interconnect_0_button_s1_readdata),             //                                                      .readdata
		.button_s1_writedata                                         (mm_interconnect_0_button_s1_writedata),            //                                                      .writedata
		.button_s1_chipselect                                        (mm_interconnect_0_button_s1_chipselect),           //                                                      .chipselect
		.bypass_sel_s1_address                                       (mm_interconnect_0_bypass_sel_s1_address),          //                                         bypass_sel_s1.address
		.bypass_sel_s1_write                                         (mm_interconnect_0_bypass_sel_s1_write),            //                                                      .write
		.bypass_sel_s1_readdata                                      (mm_interconnect_0_bypass_sel_s1_readdata),         //                                                      .readdata
		.bypass_sel_s1_writedata                                     (mm_interconnect_0_bypass_sel_s1_writedata),        //                                                      .writedata
		.bypass_sel_s1_chipselect                                    (mm_interconnect_0_bypass_sel_s1_chipselect),       //                                                      .chipselect
		.delay_lenght_s1_address                                     (mm_interconnect_0_delay_lenght_s1_address),        //                                       delay_lenght_s1.address
		.delay_lenght_s1_write                                       (mm_interconnect_0_delay_lenght_s1_write),          //                                                      .write
		.delay_lenght_s1_readdata                                    (mm_interconnect_0_delay_lenght_s1_readdata),       //                                                      .readdata
		.delay_lenght_s1_writedata                                   (mm_interconnect_0_delay_lenght_s1_writedata),      //                                                      .writedata
		.delay_lenght_s1_chipselect                                  (mm_interconnect_0_delay_lenght_s1_chipselect),     //                                                      .chipselect
		.DownSampleMult_s1_address                                   (mm_interconnect_0_downsamplemult_s1_address),      //                                     DownSampleMult_s1.address
		.DownSampleMult_s1_write                                     (mm_interconnect_0_downsamplemult_s1_write),        //                                                      .write
		.DownSampleMult_s1_readdata                                  (mm_interconnect_0_downsamplemult_s1_readdata),     //                                                      .readdata
		.DownSampleMult_s1_writedata                                 (mm_interconnect_0_downsamplemult_s1_writedata),    //                                                      .writedata
		.DownSampleMult_s1_chipselect                                (mm_interconnect_0_downsamplemult_s1_chipselect),   //                                                      .chipselect
		.fifo_memory_in_write                                        (mm_interconnect_0_fifo_memory_in_write),           //                                        fifo_memory_in.write
		.fifo_memory_in_writedata                                    (mm_interconnect_0_fifo_memory_in_writedata),       //                                                      .writedata
		.fifo_memory_in_waitrequest                                  (mm_interconnect_0_fifo_memory_in_waitrequest),     //                                                      .waitrequest
		.fifo_memory_in_csr_address                                  (mm_interconnect_0_fifo_memory_in_csr_address),     //                                    fifo_memory_in_csr.address
		.fifo_memory_in_csr_write                                    (mm_interconnect_0_fifo_memory_in_csr_write),       //                                                      .write
		.fifo_memory_in_csr_read                                     (mm_interconnect_0_fifo_memory_in_csr_read),        //                                                      .read
		.fifo_memory_in_csr_readdata                                 (mm_interconnect_0_fifo_memory_in_csr_readdata),    //                                                      .readdata
		.fifo_memory_in_csr_writedata                                (mm_interconnect_0_fifo_memory_in_csr_writedata),   //                                                      .writedata
		.fifo_memory_out_read                                        (mm_interconnect_0_fifo_memory_out_read),           //                                       fifo_memory_out.read
		.fifo_memory_out_readdata                                    (mm_interconnect_0_fifo_memory_out_readdata),       //                                                      .readdata
		.fifo_memory_out_waitrequest                                 (mm_interconnect_0_fifo_memory_out_waitrequest),    //                                                      .waitrequest
		.fir_memory_s1_address                                       (mm_interconnect_0_fir_memory_s1_address),          //                                         fir_memory_s1.address
		.fir_memory_s1_write                                         (mm_interconnect_0_fir_memory_s1_write),            //                                                      .write
		.fir_memory_s1_readdata                                      (mm_interconnect_0_fir_memory_s1_readdata),         //                                                      .readdata
		.fir_memory_s1_writedata                                     (mm_interconnect_0_fir_memory_s1_writedata),        //                                                      .writedata
		.fir_memory_s1_byteenable                                    (mm_interconnect_0_fir_memory_s1_byteenable),       //                                                      .byteenable
		.fir_memory_s1_chipselect                                    (mm_interconnect_0_fir_memory_s1_chipselect),       //                                                      .chipselect
		.fir_memory_s1_clken                                         (mm_interconnect_0_fir_memory_s1_clken),            //                                                      .clken
		.Interpo_4_0_s1_address                                      (mm_interconnect_0_interpo_4_0_s1_address),         //                                        Interpo_4_0_s1.address
		.Interpo_4_0_s1_write                                        (mm_interconnect_0_interpo_4_0_s1_write),           //                                                      .write
		.Interpo_4_0_s1_readdata                                     (mm_interconnect_0_interpo_4_0_s1_readdata),        //                                                      .readdata
		.Interpo_4_0_s1_writedata                                    (mm_interconnect_0_interpo_4_0_s1_writedata),       //                                                      .writedata
		.Interpo_4_0_s1_byteenable                                   (mm_interconnect_0_interpo_4_0_s1_byteenable),      //                                                      .byteenable
		.Interpo_4_0_s1_chipselect                                   (mm_interconnect_0_interpo_4_0_s1_chipselect),      //                                                      .chipselect
		.Interpo_4_0_s1_clken                                        (mm_interconnect_0_interpo_4_0_s1_clken),           //                                                      .clken
		.Interpo_5_0_s1_address                                      (mm_interconnect_0_interpo_5_0_s1_address),         //                                        Interpo_5_0_s1.address
		.Interpo_5_0_s1_write                                        (mm_interconnect_0_interpo_5_0_s1_write),           //                                                      .write
		.Interpo_5_0_s1_readdata                                     (mm_interconnect_0_interpo_5_0_s1_readdata),        //                                                      .readdata
		.Interpo_5_0_s1_writedata                                    (mm_interconnect_0_interpo_5_0_s1_writedata),       //                                                      .writedata
		.Interpo_5_0_s1_byteenable                                   (mm_interconnect_0_interpo_5_0_s1_byteenable),      //                                                      .byteenable
		.Interpo_5_0_s1_chipselect                                   (mm_interconnect_0_interpo_5_0_s1_chipselect),      //                                                      .chipselect
		.Interpo_5_0_s1_clken                                        (mm_interconnect_0_interpo_5_0_s1_clken),           //                                                      .clken
		.Interpo_5_1_s1_address                                      (mm_interconnect_0_interpo_5_1_s1_address),         //                                        Interpo_5_1_s1.address
		.Interpo_5_1_s1_write                                        (mm_interconnect_0_interpo_5_1_s1_write),           //                                                      .write
		.Interpo_5_1_s1_readdata                                     (mm_interconnect_0_interpo_5_1_s1_readdata),        //                                                      .readdata
		.Interpo_5_1_s1_writedata                                    (mm_interconnect_0_interpo_5_1_s1_writedata),       //                                                      .writedata
		.Interpo_5_1_s1_byteenable                                   (mm_interconnect_0_interpo_5_1_s1_byteenable),      //                                                      .byteenable
		.Interpo_5_1_s1_chipselect                                   (mm_interconnect_0_interpo_5_1_s1_chipselect),      //                                                      .chipselect
		.Interpo_5_1_s1_clken                                        (mm_interconnect_0_interpo_5_1_s1_clken),           //                                                      .clken
		.Interpo_5_2_s1_address                                      (mm_interconnect_0_interpo_5_2_s1_address),         //                                        Interpo_5_2_s1.address
		.Interpo_5_2_s1_write                                        (mm_interconnect_0_interpo_5_2_s1_write),           //                                                      .write
		.Interpo_5_2_s1_readdata                                     (mm_interconnect_0_interpo_5_2_s1_readdata),        //                                                      .readdata
		.Interpo_5_2_s1_writedata                                    (mm_interconnect_0_interpo_5_2_s1_writedata),       //                                                      .writedata
		.Interpo_5_2_s1_byteenable                                   (mm_interconnect_0_interpo_5_2_s1_byteenable),      //                                                      .byteenable
		.Interpo_5_2_s1_chipselect                                   (mm_interconnect_0_interpo_5_2_s1_chipselect),      //                                                      .chipselect
		.Interpo_5_2_s1_clken                                        (mm_interconnect_0_interpo_5_2_s1_clken),           //                                                      .clken
		.Interpo_5_3_s1_address                                      (mm_interconnect_0_interpo_5_3_s1_address),         //                                        Interpo_5_3_s1.address
		.Interpo_5_3_s1_write                                        (mm_interconnect_0_interpo_5_3_s1_write),           //                                                      .write
		.Interpo_5_3_s1_readdata                                     (mm_interconnect_0_interpo_5_3_s1_readdata),        //                                                      .readdata
		.Interpo_5_3_s1_writedata                                    (mm_interconnect_0_interpo_5_3_s1_writedata),       //                                                      .writedata
		.Interpo_5_3_s1_byteenable                                   (mm_interconnect_0_interpo_5_3_s1_byteenable),      //                                                      .byteenable
		.Interpo_5_3_s1_chipselect                                   (mm_interconnect_0_interpo_5_3_s1_chipselect),      //                                                      .chipselect
		.Interpo_5_3_s1_clken                                        (mm_interconnect_0_interpo_5_3_s1_clken),           //                                                      .clken
		.led_s1_address                                              (mm_interconnect_0_led_s1_address),                 //                                                led_s1.address
		.led_s1_write                                                (mm_interconnect_0_led_s1_write),                   //                                                      .write
		.led_s1_readdata                                             (mm_interconnect_0_led_s1_readdata),                //                                                      .readdata
		.led_s1_writedata                                            (mm_interconnect_0_led_s1_writedata),               //                                                      .writedata
		.led_s1_chipselect                                           (mm_interconnect_0_led_s1_chipselect),              //                                                      .chipselect
		.micFilter_adjust_s1_address                                 (mm_interconnect_0_micfilter_adjust_s1_address),    //                                   micFilter_adjust_s1.address
		.micFilter_adjust_s1_write                                   (mm_interconnect_0_micfilter_adjust_s1_write),      //                                                      .write
		.micFilter_adjust_s1_readdata                                (mm_interconnect_0_micfilter_adjust_s1_readdata),   //                                                      .readdata
		.micFilter_adjust_s1_writedata                               (mm_interconnect_0_micfilter_adjust_s1_writedata),  //                                                      .writedata
		.micFilter_adjust_s1_chipselect                              (mm_interconnect_0_micfilter_adjust_s1_chipselect), //                                                      .chipselect
		.micFilter_cntl_s1_address                                   (mm_interconnect_0_micfilter_cntl_s1_address),      //                                     micFilter_cntl_s1.address
		.micFilter_cntl_s1_write                                     (mm_interconnect_0_micfilter_cntl_s1_write),        //                                                      .write
		.micFilter_cntl_s1_readdata                                  (mm_interconnect_0_micfilter_cntl_s1_readdata),     //                                                      .readdata
		.micFilter_cntl_s1_writedata                                 (mm_interconnect_0_micfilter_cntl_s1_writedata),    //                                                      .writedata
		.micFilter_cntl_s1_chipselect                                (mm_interconnect_0_micfilter_cntl_s1_chipselect),   //                                                      .chipselect
		.micFilter_rst_s1_address                                    (mm_interconnect_0_micfilter_rst_s1_address),       //                                      micFilter_rst_s1.address
		.micFilter_rst_s1_write                                      (mm_interconnect_0_micfilter_rst_s1_write),         //                                                      .write
		.micFilter_rst_s1_readdata                                   (mm_interconnect_0_micfilter_rst_s1_readdata),      //                                                      .readdata
		.micFilter_rst_s1_writedata                                  (mm_interconnect_0_micfilter_rst_s1_writedata),     //                                                      .writedata
		.micFilter_rst_s1_chipselect                                 (mm_interconnect_0_micfilter_rst_s1_chipselect),    //                                                      .chipselect
		.output1_sel_s1_address                                      (mm_interconnect_0_output1_sel_s1_address),         //                                        output1_sel_s1.address
		.output1_sel_s1_write                                        (mm_interconnect_0_output1_sel_s1_write),           //                                                      .write
		.output1_sel_s1_readdata                                     (mm_interconnect_0_output1_sel_s1_readdata),        //                                                      .readdata
		.output1_sel_s1_writedata                                    (mm_interconnect_0_output1_sel_s1_writedata),       //                                                      .writedata
		.output1_sel_s1_chipselect                                   (mm_interconnect_0_output1_sel_s1_chipselect),      //                                                      .chipselect
		.output2_sel_s1_address                                      (mm_interconnect_0_output2_sel_s1_address),         //                                        output2_sel_s1.address
		.output2_sel_s1_write                                        (mm_interconnect_0_output2_sel_s1_write),           //                                                      .write
		.output2_sel_s1_readdata                                     (mm_interconnect_0_output2_sel_s1_readdata),        //                                                      .readdata
		.output2_sel_s1_writedata                                    (mm_interconnect_0_output2_sel_s1_writedata),       //                                                      .writedata
		.output2_sel_s1_chipselect                                   (mm_interconnect_0_output2_sel_s1_chipselect),      //                                                      .chipselect
		.pcie_ip_txs_address                                         (mm_interconnect_0_pcie_ip_txs_address),            //                                           pcie_ip_txs.address
		.pcie_ip_txs_write                                           (mm_interconnect_0_pcie_ip_txs_write),              //                                                      .write
		.pcie_ip_txs_read                                            (mm_interconnect_0_pcie_ip_txs_read),               //                                                      .read
		.pcie_ip_txs_readdata                                        (mm_interconnect_0_pcie_ip_txs_readdata),           //                                                      .readdata
		.pcie_ip_txs_writedata                                       (mm_interconnect_0_pcie_ip_txs_writedata),          //                                                      .writedata
		.pcie_ip_txs_burstcount                                      (mm_interconnect_0_pcie_ip_txs_burstcount),         //                                                      .burstcount
		.pcie_ip_txs_byteenable                                      (mm_interconnect_0_pcie_ip_txs_byteenable),         //                                                      .byteenable
		.pcie_ip_txs_readdatavalid                                   (mm_interconnect_0_pcie_ip_txs_readdatavalid),      //                                                      .readdatavalid
		.pcie_ip_txs_waitrequest                                     (mm_interconnect_0_pcie_ip_txs_waitrequest),        //                                                      .waitrequest
		.pcie_ip_txs_chipselect                                      (mm_interconnect_0_pcie_ip_txs_chipselect),         //                                                      .chipselect
		.sub_factor_s1_address                                       (mm_interconnect_0_sub_factor_s1_address),          //                                         sub_factor_s1.address
		.sub_factor_s1_write                                         (mm_interconnect_0_sub_factor_s1_write),            //                                                      .write
		.sub_factor_s1_readdata                                      (mm_interconnect_0_sub_factor_s1_readdata),         //                                                      .readdata
		.sub_factor_s1_writedata                                     (mm_interconnect_0_sub_factor_s1_writedata),        //                                                      .writedata
		.sub_factor_s1_chipselect                                    (mm_interconnect_0_sub_factor_s1_chipselect)        //                                                      .chipselect
	);

	de2i_150_qsys_mm_interconnect_1 mm_interconnect_1 (
		.pcie_ip_pcie_core_clk_clk                                 (pcie_ip_pcie_core_clk_clk),                 //                               pcie_ip_pcie_core_clk.clk
		.pcie_ip_bar2_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),        // pcie_ip_bar2_translator_reset_reset_bridge_in_reset.reset
		.sgdma_reset_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),            //                   sgdma_reset_reset_bridge_in_reset.reset
		.pcie_ip_bar2_address                                      (pcie_ip_bar2_address),                      //                                        pcie_ip_bar2.address
		.pcie_ip_bar2_waitrequest                                  (pcie_ip_bar2_waitrequest),                  //                                                    .waitrequest
		.pcie_ip_bar2_burstcount                                   (pcie_ip_bar2_burstcount),                   //                                                    .burstcount
		.pcie_ip_bar2_byteenable                                   (pcie_ip_bar2_byteenable),                   //                                                    .byteenable
		.pcie_ip_bar2_read                                         (pcie_ip_bar2_read),                         //                                                    .read
		.pcie_ip_bar2_readdata                                     (pcie_ip_bar2_readdata),                     //                                                    .readdata
		.pcie_ip_bar2_readdatavalid                                (pcie_ip_bar2_readdatavalid),                //                                                    .readdatavalid
		.pcie_ip_bar2_write                                        (pcie_ip_bar2_write),                        //                                                    .write
		.pcie_ip_bar2_writedata                                    (pcie_ip_bar2_writedata),                    //                                                    .writedata
		.pcie_ip_cra_address                                       (mm_interconnect_1_pcie_ip_cra_address),     //                                         pcie_ip_cra.address
		.pcie_ip_cra_write                                         (mm_interconnect_1_pcie_ip_cra_write),       //                                                    .write
		.pcie_ip_cra_read                                          (mm_interconnect_1_pcie_ip_cra_read),        //                                                    .read
		.pcie_ip_cra_readdata                                      (mm_interconnect_1_pcie_ip_cra_readdata),    //                                                    .readdata
		.pcie_ip_cra_writedata                                     (mm_interconnect_1_pcie_ip_cra_writedata),   //                                                    .writedata
		.pcie_ip_cra_byteenable                                    (mm_interconnect_1_pcie_ip_cra_byteenable),  //                                                    .byteenable
		.pcie_ip_cra_waitrequest                                   (mm_interconnect_1_pcie_ip_cra_waitrequest), //                                                    .waitrequest
		.pcie_ip_cra_chipselect                                    (mm_interconnect_1_pcie_ip_cra_chipselect),  //                                                    .chipselect
		.sgdma_csr_address                                         (mm_interconnect_1_sgdma_csr_address),       //                                           sgdma_csr.address
		.sgdma_csr_write                                           (mm_interconnect_1_sgdma_csr_write),         //                                                    .write
		.sgdma_csr_read                                            (mm_interconnect_1_sgdma_csr_read),          //                                                    .read
		.sgdma_csr_readdata                                        (mm_interconnect_1_sgdma_csr_readdata),      //                                                    .readdata
		.sgdma_csr_writedata                                       (mm_interconnect_1_sgdma_csr_writedata),     //                                                    .writedata
		.sgdma_csr_chipselect                                      (mm_interconnect_1_sgdma_csr_chipselect)     //                                                    .chipselect
	);

	de2i_150_qsys_irq_mapper irq_mapper (
		.clk           (pcie_ip_pcie_core_clk_clk),          //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.sender_irq    (pcie_ip_rxm_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~pcie_ip_pcie_core_reset_reset),     // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.clk            (pcie_ip_pcie_core_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~pcie_ip_pcie_core_reset_reset),     // reset_in0.reset
		.clk            (pcie_ip_pcie_core_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
